module sbox(
    clk,
    t0,
    t1,
    r0,
    r1,
    r2,
    r3,
    r4,
    r5,
    r6,
    r7,
    r8,
    r9,
    r10,
    r11,
    r12,
    r13,
    r14,
    r15,
    r16,
    r17,
    r18,
    r19,
    r20,
    r21,
    r22,
    r23,
    r24,
    r25,
    r26,
    r27,
    r28,
    r29,
    r30,
    r31,
    r32,
    r33,
    r34,
    r35,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_16,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    y0,
    y1,
);
//INPUTS
    input clk;
    input  [31:0] t0;
    input  [31:0] t1;
    input  [31:0] r0;
    input  [31:0] r1;
    input  [31:0] r2;
    input  [31:0] r3;
    input  [31:0] r4;
    input  [31:0] r5;
    input  [31:0] r6;
    input  [31:0] r7;
    input  [31:0] r8;
    input  [31:0] r9;
    input  [31:0] r10;
    input  [31:0] r11;
    input  [31:0] r12;
    input  [31:0] r13;
    input  [31:0] r14;
    input  [31:0] r15;
    input  [31:0] r16;
    input  [31:0] r17;
    input  [31:0] r18;
    input  [31:0] r19;
    input  [31:0] r20;
    input  [31:0] r21;
    input  [31:0] r22;
    input  [31:0] r23;
    input  [31:0] r24;
    input  [31:0] r25;
    input  [31:0] r26;
    input  [31:0] r27;
    input  [31:0] r28;
    input  [31:0] r29;
    input  [31:0] r30;
    input  [31:0] r31;
    input  [31:0] r32;
    input  [31:0] r33;
    input  [31:0] r34;
    input  [31:0] r35;
    input  [31:0] dec_0;
    input  [31:0] dec_1;
    input  [31:0] dec_255;
    input  [31:0] dec_169;
    input  [31:0] dec_129;
    input  [31:0] dec_9;
    input  [31:0] dec_72;
    input  [31:0] dec_242;
    input  [31:0] dec_243;
    input  [31:0] dec_152;
    input  [31:0] dec_240;
    input  [31:0] dec_4;
    input  [31:0] dec_15;
    input  [31:0] dec_12;
    input  [31:0] dec_2;
    input  [31:0] dec_3;
    input  [31:0] dec_16;
    input  [31:0] dec_36;
    input  [31:0] dec_220;
    input  [31:0] dec_11;
    input  [31:0] dec_158;
    input  [31:0] dec_45;
    input  [31:0] dec_88;
    input  [31:0] dec_99;
//OUTPUTS
    output reg  [31:0] y0;
    output reg  [31:0] y1;
//Intermediate values
    wire [31:0] z2945_assgn2945;
    reg [31:0] z2945_assgn29450;
    reg [31:0] z2945_assgn29451;
    reg [31:0] z2945_assgn29452;
    reg [31:0] z2945_assgn29453;
    reg [31:0] z2945_assgn29454;
    reg [31:0] z2945_assgn29455;
    reg [31:0] z2945_assgn29456;
    reg [31:0] z2945_assgn29457;
    reg [31:0] z2945_assgn29458;
    reg [31:0] dec_99_inp;
    wire [31:0] z2947_assgn2947;
    reg [31:0] z2947_assgn29470;
    reg [31:0] z2947_assgn29471;
    reg [31:0] z2947_assgn29472;
    reg [31:0] z2947_assgn29473;
    reg [31:0] z2947_assgn29474;
    reg [31:0] z2947_assgn29475;
    reg [31:0] z2947_assgn29476;
    reg [31:0] z2947_assgn29477;
    reg [31:0] z2947_assgn29478;
    reg [31:0] dec_88_inp;
    wire [31:0] z2949_assgn2949;
    reg [31:0] z2949_assgn29490;
    reg [31:0] z2949_assgn29491;
    reg [31:0] z2949_assgn29492;
    reg [31:0] z2949_assgn29493;
    reg [31:0] z2949_assgn29494;
    reg [31:0] z2949_assgn29495;
    reg [31:0] z2949_assgn29496;
    reg [31:0] z2949_assgn29497;
    reg [31:0] z2949_assgn29498;
    reg [31:0] dec_45_inp;
    wire [31:0] z2951_assgn2951;
    reg [31:0] z2951_assgn29510;
    reg [31:0] z2951_assgn29511;
    reg [31:0] z2951_assgn29512;
    reg [31:0] z2951_assgn29513;
    reg [31:0] z2951_assgn29514;
    reg [31:0] z2951_assgn29515;
    reg [31:0] z2951_assgn29516;
    reg [31:0] z2951_assgn29517;
    reg [31:0] z2951_assgn29518;
    reg [31:0] dec_158_inp;
    wire [31:0] z2953_assgn2953;
    reg [31:0] z2953_assgn29530;
    reg [31:0] z2953_assgn29531;
    reg [31:0] z2953_assgn29532;
    reg [31:0] z2953_assgn29533;
    reg [31:0] z2953_assgn29534;
    reg [31:0] z2953_assgn29535;
    reg [31:0] z2953_assgn29536;
    reg [31:0] z2953_assgn29537;
    reg [31:0] z2953_assgn29538;
    reg [31:0] dec_11_inp;
    wire [31:0] z2955_assgn2955;
    reg [31:0] z2955_assgn29550;
    reg [31:0] z2955_assgn29551;
    reg [31:0] z2955_assgn29552;
    reg [31:0] z2955_assgn29553;
    reg [31:0] z2955_assgn29554;
    reg [31:0] z2955_assgn29555;
    reg [31:0] z2955_assgn29556;
    reg [31:0] z2955_assgn29557;
    reg [31:0] z2955_assgn29558;
    reg [31:0] dec_220_inp;
    wire [31:0] z2957_assgn2957;
    reg [31:0] z2957_assgn29570;
    reg [31:0] z2957_assgn29571;
    reg [31:0] z2957_assgn29572;
    reg [31:0] z2957_assgn29573;
    reg [31:0] z2957_assgn29574;
    reg [31:0] z2957_assgn29575;
    reg [31:0] z2957_assgn29576;
    reg [31:0] z2957_assgn29577;
    reg [31:0] z2957_assgn29578;
    reg [31:0] dec_36_inp;
    wire [31:0] dec_16_inp;
    reg [31:0] z1_assgn1;
    wire [31:0] dec_3_inp;
    wire [31:0] dec_2_inp;
    wire [31:0] dec_12_inp;
    wire [31:0] dec_15_inp;
    wire [31:0] dec_4_inp;
    reg [31:0] z3_assgn3;
    wire [31:0] z2975_assgn2975;
    reg [31:0] z2975_assgn29750;
    reg [31:0] z2975_assgn29751;
    reg [31:0] dec_240_inp;
    wire [31:0] dec_152_inp;
    wire [31:0] dec_243_inp;
    wire [31:0] dec_242_inp;
    wire [31:0] dec_72_inp;
    wire [31:0] dec_9_inp;
    wire [31:0] dec_129_inp;
    wire [31:0] dec_169_inp;
    wire [31:0] dec_255_inp;
    wire [31:0] dec_1_inp;
    wire [31:0] dec_0_inp;
    wire [31:0] t0_inp;
    wire [31:0] t1_inp;
    wire [31:0] r0_inp;
    reg [31:0] z5_assgn5;
    wire [31:0] r1_inp;
    reg [31:0] z7_assgn7;
    wire [31:0] r2_inp;
    reg [31:0] z9_assgn9;
    wire [31:0] r3_inp;
    reg [31:0] z11_assgn11;
    wire [31:0] r4_inp;
    reg [31:0] z13_assgn13;
    wire [31:0] r5_inp;
    reg [31:0] z15_assgn15;
    wire [31:0] r6_inp;
    reg [31:0] z17_assgn17;
    wire [31:0] r7_inp;
    reg [31:0] z19_assgn19;
    wire [31:0] r8_inp;
    reg [31:0] z21_assgn21;
    wire [31:0] z3037_assgn3037;
    reg [31:0] z3037_assgn30370;
    reg [31:0] z3037_assgn30371;
    reg [31:0] z3037_assgn30372;
    reg [31:0] z3037_assgn30373;
    reg [31:0] r9_inp;
    wire [31:0] z3039_assgn3039;
    reg [31:0] z3039_assgn30390;
    reg [31:0] z3039_assgn30391;
    reg [31:0] z3039_assgn30392;
    reg [31:0] z3039_assgn30393;
    reg [31:0] r10_inp;
    wire [31:0] z3041_assgn3041;
    reg [31:0] z3041_assgn30410;
    reg [31:0] z3041_assgn30411;
    reg [31:0] z3041_assgn30412;
    reg [31:0] z3041_assgn30413;
    reg [31:0] r11_inp;
    wire [31:0] z3043_assgn3043;
    reg [31:0] z3043_assgn30430;
    reg [31:0] z3043_assgn30431;
    reg [31:0] z3043_assgn30432;
    reg [31:0] z3043_assgn30433;
    reg [31:0] z3043_assgn30434;
    reg [31:0] r12_inp;
    wire [31:0] z3045_assgn3045;
    reg [31:0] z3045_assgn30450;
    reg [31:0] z3045_assgn30451;
    reg [31:0] z3045_assgn30452;
    reg [31:0] z3045_assgn30453;
    reg [31:0] z3045_assgn30454;
    reg [31:0] r13_inp;
    wire [31:0] z3047_assgn3047;
    reg [31:0] z3047_assgn30470;
    reg [31:0] z3047_assgn30471;
    reg [31:0] z3047_assgn30472;
    reg [31:0] z3047_assgn30473;
    reg [31:0] z3047_assgn30474;
    reg [31:0] r14_inp;
    wire [31:0] z3049_assgn3049;
    reg [31:0] z3049_assgn30490;
    reg [31:0] z3049_assgn30491;
    reg [31:0] z3049_assgn30492;
    reg [31:0] z3049_assgn30493;
    reg [31:0] z3049_assgn30494;
    reg [31:0] r15_inp;
    wire [31:0] z3051_assgn3051;
    reg [31:0] z3051_assgn30510;
    reg [31:0] z3051_assgn30511;
    reg [31:0] z3051_assgn30512;
    reg [31:0] z3051_assgn30513;
    reg [31:0] z3051_assgn30514;
    reg [31:0] r16_inp;
    wire [31:0] z3053_assgn3053;
    reg [31:0] z3053_assgn30530;
    reg [31:0] z3053_assgn30531;
    reg [31:0] z3053_assgn30532;
    reg [31:0] z3053_assgn30533;
    reg [31:0] z3053_assgn30534;
    reg [31:0] r17_inp;
    wire [31:0] z3055_assgn3055;
    reg [31:0] z3055_assgn30550;
    reg [31:0] z3055_assgn30551;
    reg [31:0] z3055_assgn30552;
    reg [31:0] z3055_assgn30553;
    reg [31:0] z3055_assgn30554;
    reg [31:0] z3055_assgn30555;
    reg [31:0] r18_inp;
    wire [31:0] z3057_assgn3057;
    reg [31:0] z3057_assgn30570;
    reg [31:0] z3057_assgn30571;
    reg [31:0] z3057_assgn30572;
    reg [31:0] z3057_assgn30573;
    reg [31:0] z3057_assgn30574;
    reg [31:0] z3057_assgn30575;
    reg [31:0] r19_inp;
    wire [31:0] z3059_assgn3059;
    reg [31:0] z3059_assgn30590;
    reg [31:0] z3059_assgn30591;
    reg [31:0] z3059_assgn30592;
    reg [31:0] z3059_assgn30593;
    reg [31:0] z3059_assgn30594;
    reg [31:0] z3059_assgn30595;
    reg [31:0] r20_inp;
    wire [31:0] z3061_assgn3061;
    reg [31:0] z3061_assgn30610;
    reg [31:0] z3061_assgn30611;
    reg [31:0] z3061_assgn30612;
    reg [31:0] z3061_assgn30613;
    reg [31:0] z3061_assgn30614;
    reg [31:0] z3061_assgn30615;
    reg [31:0] r21_inp;
    wire [31:0] z3063_assgn3063;
    reg [31:0] z3063_assgn30630;
    reg [31:0] z3063_assgn30631;
    reg [31:0] z3063_assgn30632;
    reg [31:0] z3063_assgn30633;
    reg [31:0] z3063_assgn30634;
    reg [31:0] z3063_assgn30635;
    reg [31:0] r22_inp;
    wire [31:0] z3065_assgn3065;
    reg [31:0] z3065_assgn30650;
    reg [31:0] z3065_assgn30651;
    reg [31:0] z3065_assgn30652;
    reg [31:0] z3065_assgn30653;
    reg [31:0] z3065_assgn30654;
    reg [31:0] z3065_assgn30655;
    reg [31:0] r23_inp;
    wire [31:0] z3067_assgn3067;
    reg [31:0] z3067_assgn30670;
    reg [31:0] z3067_assgn30671;
    reg [31:0] z3067_assgn30672;
    reg [31:0] z3067_assgn30673;
    reg [31:0] z3067_assgn30674;
    reg [31:0] z3067_assgn30675;
    reg [31:0] r24_inp;
    wire [31:0] z3069_assgn3069;
    reg [31:0] z3069_assgn30690;
    reg [31:0] z3069_assgn30691;
    reg [31:0] z3069_assgn30692;
    reg [31:0] z3069_assgn30693;
    reg [31:0] z3069_assgn30694;
    reg [31:0] z3069_assgn30695;
    reg [31:0] r25_inp;
    wire [31:0] z3071_assgn3071;
    reg [31:0] z3071_assgn30710;
    reg [31:0] z3071_assgn30711;
    reg [31:0] z3071_assgn30712;
    reg [31:0] z3071_assgn30713;
    reg [31:0] z3071_assgn30714;
    reg [31:0] z3071_assgn30715;
    reg [31:0] r26_inp;
    wire [31:0] z3073_assgn3073;
    reg [31:0] z3073_assgn30730;
    reg [31:0] z3073_assgn30731;
    reg [31:0] z3073_assgn30732;
    reg [31:0] z3073_assgn30733;
    reg [31:0] z3073_assgn30734;
    reg [31:0] z3073_assgn30735;
    reg [31:0] r27_inp;
    wire [31:0] z3075_assgn3075;
    reg [31:0] z3075_assgn30750;
    reg [31:0] z3075_assgn30751;
    reg [31:0] z3075_assgn30752;
    reg [31:0] z3075_assgn30753;
    reg [31:0] z3075_assgn30754;
    reg [31:0] z3075_assgn30755;
    reg [31:0] r28_inp;
    wire [31:0] z3077_assgn3077;
    reg [31:0] z3077_assgn30770;
    reg [31:0] z3077_assgn30771;
    reg [31:0] z3077_assgn30772;
    reg [31:0] z3077_assgn30773;
    reg [31:0] z3077_assgn30774;
    reg [31:0] z3077_assgn30775;
    reg [31:0] r29_inp;
    wire [31:0] z3079_assgn3079;
    reg [31:0] z3079_assgn30790;
    reg [31:0] z3079_assgn30791;
    reg [31:0] z3079_assgn30792;
    reg [31:0] z3079_assgn30793;
    reg [31:0] z3079_assgn30794;
    reg [31:0] z3079_assgn30795;
    reg [31:0] r30_inp;
    wire [31:0] z3081_assgn3081;
    reg [31:0] z3081_assgn30810;
    reg [31:0] z3081_assgn30811;
    reg [31:0] z3081_assgn30812;
    reg [31:0] z3081_assgn30813;
    reg [31:0] z3081_assgn30814;
    reg [31:0] z3081_assgn30815;
    reg [31:0] r31_inp;
    wire [31:0] z3083_assgn3083;
    reg [31:0] z3083_assgn30830;
    reg [31:0] z3083_assgn30831;
    reg [31:0] z3083_assgn30832;
    reg [31:0] z3083_assgn30833;
    reg [31:0] z3083_assgn30834;
    reg [31:0] z3083_assgn30835;
    reg [31:0] r32_inp;
    wire [31:0] z3085_assgn3085;
    reg [31:0] z3085_assgn30850;
    reg [31:0] z3085_assgn30851;
    reg [31:0] z3085_assgn30852;
    reg [31:0] z3085_assgn30853;
    reg [31:0] z3085_assgn30854;
    reg [31:0] z3085_assgn30855;
    reg [31:0] r33_inp;
    wire [31:0] z3087_assgn3087;
    reg [31:0] z3087_assgn30870;
    reg [31:0] z3087_assgn30871;
    reg [31:0] z3087_assgn30872;
    reg [31:0] z3087_assgn30873;
    reg [31:0] z3087_assgn30874;
    reg [31:0] z3087_assgn30875;
    reg [31:0] r34_inp;
    wire [31:0] z3089_assgn3089;
    reg [31:0] z3089_assgn30890;
    reg [31:0] z3089_assgn30891;
    reg [31:0] z3089_assgn30892;
    reg [31:0] z3089_assgn30893;
    reg [31:0] z3089_assgn30894;
    reg [31:0] z3089_assgn30895;
    reg [31:0] r35_inp;
    wire [31:0] y_G256_newbasis0;
    wire [31:0] tempy1_G256_newbasis0;
    wire [31:0] cond1_G256_newbasis0;
    wire [31:0] negCond1_G256_newbasis0;
    wire [31:0] yxorb1_G256_newbasis0;
    wire [31:0] ny1_G256_newbasis0;
    wire [31:0] tempyIntoNegCond1_G256_newbasis0;
    wire [31:0] y1_G256_newbasis0;
    wire [31:0] x1_G256_newbasis0;
    wire [31:0] tempy2_G256_newbasis0;
    wire [31:0] cond2_G256_newbasis0;
    wire [31:0] negCond2_G256_newbasis0;
    wire [31:0] yxorb2_G256_newbasis0;
    wire [31:0] ny2_G256_newbasis0;
    wire [31:0] tempyIntoNegCond2_G256_newbasis0;
    wire [31:0] y2_G256_newbasis0;
    wire [31:0] x2_G256_newbasis0;
    wire [31:0] tempy3_G256_newbasis0;
    wire [31:0] cond3_G256_newbasis0;
    wire [31:0] negCond3_G256_newbasis0;
    wire [31:0] yxorb3_G256_newbasis0;
    wire [31:0] ny3_G256_newbasis0;
    wire [31:0] tempyIntoNegCond3_G256_newbasis0;
    wire [31:0] y3_G256_newbasis0;
    wire [31:0] x3_G256_newbasis0;
    wire [31:0] tempy4_G256_newbasis0;
    wire [31:0] cond4_G256_newbasis0;
    wire [31:0] negCond4_G256_newbasis0;
    wire [31:0] yxorb4_G256_newbasis0;
    wire [31:0] ny4_G256_newbasis0;
    wire [31:0] tempyIntoNegCond4_G256_newbasis0;
    wire [31:0] y4_G256_newbasis0;
    wire [31:0] x4_G256_newbasis0;
    wire [31:0] tempy5_G256_newbasis0;
    wire [31:0] cond5_G256_newbasis0;
    wire [31:0] negCond5_G256_newbasis0;
    wire [31:0] yxorb5_G256_newbasis0;
    wire [31:0] ny5_G256_newbasis0;
    wire [31:0] tempyIntoNegCond5_G256_newbasis0;
    wire [31:0] y5_G256_newbasis0;
    wire [31:0] x5_G256_newbasis0;
    wire [31:0] tempy6_G256_newbasis0;
    wire [31:0] cond6_G256_newbasis0;
    wire [31:0] negCond6_G256_newbasis0;
    wire [31:0] yxorb6_G256_newbasis0;
    wire [31:0] ny6_G256_newbasis0;
    wire [31:0] tempyIntoNegCond6_G256_newbasis0;
    wire [31:0] y6_G256_newbasis0;
    wire [31:0] x6_G256_newbasis0;
    wire [31:0] tempy7_G256_newbasis0;
    wire [31:0] cond7_G256_newbasis0;
    wire [31:0] negCond7_G256_newbasis0;
    wire [31:0] yxorb7_G256_newbasis0;
    wire [31:0] ny7_G256_newbasis0;
    wire [31:0] tempyIntoNegCond7_G256_newbasis0;
    wire [31:0] y7_G256_newbasis0;
    wire [31:0] x7_G256_newbasis0;
    wire [31:0] tempy8_G256_newbasis0;
    wire [31:0] cond8_G256_newbasis0;
    wire [31:0] negCond8_G256_newbasis0;
    wire [31:0] yxorb8_G256_newbasis0;
    wire [31:0] ny8_G256_newbasis0;
    wire [31:0] tempyIntoNegCond8_G256_newbasis0;
    wire [31:0] y8_G256_newbasis0;
    wire [31:0] z3219_assgn3219;
    reg [31:0] z3219_assgn32190;
    reg [31:0] z3219_assgn32191;
    reg [31:0] z3219_assgn32192;
    reg [31:0] z3219_assgn32193;
    reg [31:0] z3219_assgn32194;
    reg [31:0] z3219_assgn32195;
    reg [31:0] z3219_assgn32196;
    reg [31:0] z3219_assgn32197;
    reg [31:0] z3219_assgn32198;
    reg [31:0] z297_assgn297;
    wire [31:0] z3221_assgn3221;
    reg [31:0] z3221_assgn32210;
    reg [31:0] z3221_assgn32211;
    reg [31:0] z3221_assgn32212;
    reg [31:0] z3221_assgn32213;
    reg [31:0] z3221_assgn32214;
    reg [31:0] z3221_assgn32215;
    reg [31:0] z3221_assgn32216;
    reg [31:0] z3221_assgn32217;
    reg [31:0] z3221_assgn32218;
    reg [31:0] z298_assgn298;
    wire [31:0] x8_G256_newbasis0;
    wire [31:0] t2;
    wire [31:0] z_y_G256_newbasis0;
    wire [31:0] z_tempy1_G256_newbasis0;
    wire [31:0] z_cond1_G256_newbasis0;
    wire [31:0] z_negCond1_G256_newbasis0;
    wire [31:0] z_yxorb1_G256_newbasis0;
    wire [31:0] z_ny1_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond1_G256_newbasis0;
    wire [31:0] z_y1_G256_newbasis0;
    wire [31:0] z_x1_G256_newbasis0;
    wire [31:0] z_tempy2_G256_newbasis0;
    wire [31:0] z_cond2_G256_newbasis0;
    wire [31:0] z_negCond2_G256_newbasis0;
    wire [31:0] z_yxorb2_G256_newbasis0;
    wire [31:0] z_ny2_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond2_G256_newbasis0;
    wire [31:0] z_y2_G256_newbasis0;
    wire [31:0] z_x2_G256_newbasis0;
    wire [31:0] z_tempy3_G256_newbasis0;
    wire [31:0] z_cond3_G256_newbasis0;
    wire [31:0] z_negCond3_G256_newbasis0;
    wire [31:0] z_yxorb3_G256_newbasis0;
    wire [31:0] z_ny3_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond3_G256_newbasis0;
    wire [31:0] z_y3_G256_newbasis0;
    wire [31:0] z_x3_G256_newbasis0;
    wire [31:0] z_tempy4_G256_newbasis0;
    wire [31:0] z_cond4_G256_newbasis0;
    wire [31:0] z_negCond4_G256_newbasis0;
    wire [31:0] z_yxorb4_G256_newbasis0;
    wire [31:0] z_ny4_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond4_G256_newbasis0;
    wire [31:0] z_y4_G256_newbasis0;
    wire [31:0] z_x4_G256_newbasis0;
    wire [31:0] z_tempy5_G256_newbasis0;
    wire [31:0] z_cond5_G256_newbasis0;
    wire [31:0] z_negCond5_G256_newbasis0;
    wire [31:0] z_yxorb5_G256_newbasis0;
    wire [31:0] z_ny5_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond5_G256_newbasis0;
    wire [31:0] z_y5_G256_newbasis0;
    wire [31:0] z_x5_G256_newbasis0;
    wire [31:0] z_tempy6_G256_newbasis0;
    wire [31:0] z_cond6_G256_newbasis0;
    wire [31:0] z_negCond6_G256_newbasis0;
    wire [31:0] z_yxorb6_G256_newbasis0;
    wire [31:0] z_ny6_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond6_G256_newbasis0;
    wire [31:0] z_y6_G256_newbasis0;
    wire [31:0] z_x6_G256_newbasis0;
    wire [31:0] z_tempy7_G256_newbasis0;
    wire [31:0] z_cond7_G256_newbasis0;
    wire [31:0] z_negCond7_G256_newbasis0;
    wire [31:0] z_yxorb7_G256_newbasis0;
    wire [31:0] z_ny7_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond7_G256_newbasis0;
    wire [31:0] z_y7_G256_newbasis0;
    wire [31:0] z_x7_G256_newbasis0;
    wire [31:0] z_tempy8_G256_newbasis0;
    wire [31:0] z_cond8_G256_newbasis0;
    wire [31:0] z_negCond8_G256_newbasis0;
    wire [31:0] z_yxorb8_G256_newbasis0;
    wire [31:0] z_ny8_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond8_G256_newbasis0;
    wire [31:0] z_y8_G256_newbasis0;
    wire [31:0] z3355_assgn3355;
    reg [31:0] z3355_assgn33550;
    reg [31:0] z3355_assgn33551;
    reg [31:0] z3355_assgn33552;
    reg [31:0] z3355_assgn33553;
    reg [31:0] z3355_assgn33554;
    reg [31:0] z3355_assgn33555;
    reg [31:0] z3355_assgn33556;
    reg [31:0] z3355_assgn33557;
    reg [31:0] z3355_assgn33558;
    reg [31:0] z429_assgn429;
    wire [31:0] z3357_assgn3357;
    reg [31:0] z3357_assgn33570;
    reg [31:0] z3357_assgn33571;
    reg [31:0] z3357_assgn33572;
    reg [31:0] z3357_assgn33573;
    reg [31:0] z3357_assgn33574;
    reg [31:0] z3357_assgn33575;
    reg [31:0] z3357_assgn33576;
    reg [31:0] z3357_assgn33577;
    reg [31:0] z3357_assgn33578;
    reg [31:0] z430_assgn430;
    wire [31:0] z_x8_G256_newbasis0;
    wire [31:0] t3;
    wire [31:0] z3363_assgn3363;
    reg [31:0] z3363_assgn33630;
    reg [31:0] z3363_assgn33631;
    reg [31:0] z434_assgn434;
    wire [31:0] a0_0_G256_inv0;
    wire [31:0] z3367_assgn3367;
    reg [31:0] z3367_assgn33670;
    reg [31:0] z3367_assgn33671;
    reg [31:0] z436_assgn436;
    wire [31:0] a1_0_G256_inv0;
    wire [31:0] z3371_assgn3371;
    reg [31:0] z3371_assgn33710;
    reg [31:0] z437_assgn437;
    wire [31:0] a0_G256_inv0;
    wire [31:0] z3375_assgn3375;
    reg [31:0] z3375_assgn33750;
    reg [31:0] z439_assgn439;
    wire [31:0] a1_G256_inv0;
    wire [31:0] b0_G256_inv0;
    wire [31:0] b1_G256_inv0;
    wire [31:0] z3383_assgn3383;
    reg [31:0] z3383_assgn33830;
    reg [31:0] z3383_assgn33831;
    reg [31:0] z3383_assgn33832;
    reg [31:0] z445_assgn445;
    reg [31:0] a0_G256_inv0_reg;
    wire [31:0] a0xorb0_G256_inv0;
    wire [31:0] z3387_assgn3387;
    reg [31:0] z3387_assgn33870;
    reg [31:0] z3387_assgn33871;
    reg [31:0] z3387_assgn33872;
    reg [31:0] z447_assgn447;
    reg [31:0] a1_G256_inv0_reg;
    wire [31:0] a1xorb1_G256_inv0;
    wire [31:0] z3391_assgn3391;
    reg [31:0] z3391_assgn33910;
    reg [31:0] z3391_assgn33911;
    reg [31:0] z3391_assgn33912;
    reg [31:0] z449_assgn449;
    wire [31:0] a0_0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3395_assgn3395;
    reg [31:0] z3395_assgn33950;
    reg [31:0] z3395_assgn33951;
    reg [31:0] z3395_assgn33952;
    reg [31:0] z451_assgn451;
    wire [31:0] a1_0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3399_assgn3399;
    reg [31:0] z3399_assgn33990;
    reg [31:0] z3399_assgn33991;
    reg [31:0] z3399_assgn33992;
    reg [31:0] z453_assgn453;
    wire [31:0] a0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3403_assgn3403;
    reg [31:0] z3403_assgn34030;
    reg [31:0] z3403_assgn34031;
    reg [31:0] z3403_assgn34032;
    reg [31:0] z455_assgn455;
    wire [31:0] a1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3407_assgn3407;
    reg [31:0] z3407_assgn34070;
    reg [31:0] z3407_assgn34071;
    reg [31:0] z3407_assgn34072;
    reg [31:0] z457_assgn457;
    wire [31:0] b0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3411_assgn3411;
    reg [31:0] z3411_assgn34110;
    reg [31:0] z3411_assgn34111;
    reg [31:0] z3411_assgn34112;
    reg [31:0] z459_assgn459;
    wire [31:0] b1_G16_sq_scl0_G256_inv0;
    wire [31:0] p0_0_G16_sq_scl0_G256_inv0;
    wire [31:0] p1_0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3419_assgn3419;
    reg [31:0] z3419_assgn34190;
    reg [31:0] z3419_assgn34191;
    reg [31:0] z3419_assgn34192;
    reg [31:0] z465_assgn465;
    wire [31:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3423_assgn3423;
    reg [31:0] z3423_assgn34230;
    reg [31:0] z3423_assgn34231;
    reg [31:0] z3423_assgn34232;
    reg [31:0] z467_assgn467;
    wire [31:0] a1_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3427_assgn3427;
    reg [31:0] z3427_assgn34270;
    reg [31:0] z3427_assgn34271;
    reg [31:0] z3427_assgn34272;
    reg [31:0] z469_assgn469;
    wire [31:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3431_assgn3431;
    reg [31:0] z3431_assgn34310;
    reg [31:0] z3431_assgn34311;
    reg [31:0] z3431_assgn34312;
    reg [31:0] z471_assgn471;
    wire [31:0] a1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3435_assgn3435;
    reg [31:0] z3435_assgn34350;
    reg [31:0] z3435_assgn34351;
    reg [31:0] z3435_assgn34352;
    reg [31:0] z473_assgn473;
    wire [31:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3439_assgn3439;
    reg [31:0] z3439_assgn34390;
    reg [31:0] z3439_assgn34391;
    reg [31:0] z3439_assgn34392;
    reg [31:0] z475_assgn475;
    wire [31:0] b1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3443_assgn3443;
    reg [31:0] z3443_assgn34430;
    reg [31:0] z3443_assgn34431;
    reg [31:0] z3443_assgn34432;
    reg [31:0] z477_assgn477;
    wire [31:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3447_assgn3447;
    reg [31:0] z3447_assgn34470;
    reg [31:0] z3447_assgn34471;
    reg [31:0] z3447_assgn34472;
    reg [31:0] z479_assgn479;
    wire [31:0] b1ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] p0_G16_sq_scl0_G256_inv0;
    wire [31:0] p1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3455_assgn3455;
    reg [31:0] z3455_assgn34550;
    reg [31:0] z3455_assgn34551;
    reg [31:0] z3455_assgn34552;
    reg [31:0] z485_assgn485;
    wire [31:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3459_assgn3459;
    reg [31:0] z3459_assgn34590;
    reg [31:0] z3459_assgn34591;
    reg [31:0] z3459_assgn34592;
    reg [31:0] z487_assgn487;
    wire [31:0] a1_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3463_assgn3463;
    reg [31:0] z3463_assgn34630;
    reg [31:0] z3463_assgn34631;
    reg [31:0] z3463_assgn34632;
    reg [31:0] z489_assgn489;
    wire [31:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3467_assgn3467;
    reg [31:0] z3467_assgn34670;
    reg [31:0] z3467_assgn34671;
    reg [31:0] z3467_assgn34672;
    reg [31:0] z491_assgn491;
    wire [31:0] a1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3471_assgn3471;
    reg [31:0] z3471_assgn34710;
    reg [31:0] z3471_assgn34711;
    reg [31:0] z3471_assgn34712;
    reg [31:0] z493_assgn493;
    wire [31:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3475_assgn3475;
    reg [31:0] z3475_assgn34750;
    reg [31:0] z3475_assgn34751;
    reg [31:0] z3475_assgn34752;
    reg [31:0] z495_assgn495;
    wire [31:0] b1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3479_assgn3479;
    reg [31:0] z3479_assgn34790;
    reg [31:0] z3479_assgn34791;
    reg [31:0] z3479_assgn34792;
    reg [31:0] z497_assgn497;
    wire [31:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3483_assgn3483;
    reg [31:0] z3483_assgn34830;
    reg [31:0] z3483_assgn34831;
    reg [31:0] z3483_assgn34832;
    reg [31:0] z499_assgn499;
    wire [31:0] b1ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] q0_0_G16_sq_scl0_G256_inv0;
    wire [31:0] q1_0_G16_sq_scl0_G256_inv0;
    wire [31:0] z3491_assgn3491;
    reg [31:0] z3491_assgn34910;
    reg [31:0] z3491_assgn34911;
    reg [31:0] z3491_assgn34912;
    reg [31:0] z505_assgn505;
    wire [31:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3495_assgn3495;
    reg [31:0] z3495_assgn34950;
    reg [31:0] z3495_assgn34951;
    reg [31:0] z3495_assgn34952;
    reg [31:0] z507_assgn507;
    wire [31:0] a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3499_assgn3499;
    reg [31:0] z3499_assgn34990;
    reg [31:0] z3499_assgn34991;
    reg [31:0] z3499_assgn34992;
    reg [31:0] z509_assgn509;
    wire [31:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3503_assgn3503;
    reg [31:0] z3503_assgn35030;
    reg [31:0] z3503_assgn35031;
    reg [31:0] z3503_assgn35032;
    reg [31:0] z511_assgn511;
    wire [31:0] a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3507_assgn3507;
    reg [31:0] z3507_assgn35070;
    reg [31:0] z3507_assgn35071;
    reg [31:0] z3507_assgn35072;
    reg [31:0] z513_assgn513;
    wire [31:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3511_assgn3511;
    reg [31:0] z3511_assgn35110;
    reg [31:0] z3511_assgn35111;
    reg [31:0] z3511_assgn35112;
    reg [31:0] z515_assgn515;
    wire [31:0] b1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] p1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] q1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3523_assgn3523;
    reg [31:0] z3523_assgn35230;
    reg [31:0] z3523_assgn35231;
    reg [31:0] z3523_assgn35232;
    reg [31:0] z525_assgn525;
    wire [31:0] p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] z3527_assgn3527;
    reg [31:0] z3527_assgn35270;
    reg [31:0] z3527_assgn35271;
    reg [31:0] z3527_assgn35272;
    reg [31:0] z527_assgn527;
    wire [31:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] q0_G16_sq_scl0_G256_inv0;
    wire [31:0] q1_G16_sq_scl0_G256_inv0;
    wire [31:0] z3535_assgn3535;
    reg [31:0] z3535_assgn35350;
    reg [31:0] z3535_assgn35351;
    reg [31:0] z3535_assgn35352;
    reg [31:0] z533_assgn533;
    wire [31:0] p0ls2_G16_sq_scl0_G256_inv0;
    wire [31:0] z3539_assgn3539;
    reg [31:0] z3539_assgn35390;
    reg [31:0] z3539_assgn35391;
    reg [31:0] z3539_assgn35392;
    reg [31:0] z535_assgn535;
    wire [31:0] p1ls2_G16_sq_scl0_G256_inv0;
    wire [31:0] c0_G256_inv0;
    wire [31:0] c1_G256_inv0;
    wire [31:0] r00_G16_mul0_G256_inv0;
    wire [31:0] r10_G16_mul0_G256_inv0;
    wire [31:0] r20_G16_mul0_G256_inv0;
    wire [31:0] r30_G16_mul0_G256_inv0;
    wire [31:0] r40_G16_mul0_G256_inv0;
    wire [31:0] r50_G16_mul0_G256_inv0;
    wire [31:0] r60_G16_mul0_G256_inv0;
    wire [31:0] r70_G16_mul0_G256_inv0;
    wire [31:0] r80_G16_mul0_G256_inv0;
    wire [31:0] z3565_assgn3565;
    reg [31:0] z3565_assgn35650;
    reg [31:0] z3565_assgn35651;
    reg [31:0] z559_assgn559;
    wire [31:0] a0_0_G16_mul0_G256_inv0;
    wire [31:0] z3569_assgn3569;
    reg [31:0] z3569_assgn35690;
    reg [31:0] z3569_assgn35691;
    reg [31:0] z561_assgn561;
    wire [31:0] a1_0_G16_mul0_G256_inv0;
    wire [31:0] z3573_assgn3573;
    reg [31:0] z3573_assgn35730;
    reg [31:0] z3573_assgn35731;
    reg [31:0] z563_assgn563;
    wire [31:0] a0_G16_mul0_G256_inv0;
    wire [31:0] z3577_assgn3577;
    reg [31:0] z3577_assgn35770;
    reg [31:0] z3577_assgn35771;
    reg [31:0] z565_assgn565;
    wire [31:0] a1_G16_mul0_G256_inv0;
    wire [31:0] z3581_assgn3581;
    reg [31:0] z3581_assgn35810;
    reg [31:0] z3581_assgn35811;
    reg [31:0] z567_assgn567;
    wire [31:0] b0_G16_mul0_G256_inv0;
    wire [31:0] z3585_assgn3585;
    reg [31:0] z3585_assgn35850;
    reg [31:0] z3585_assgn35851;
    reg [31:0] z569_assgn569;
    wire [31:0] b1_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G16_mul0_G256_inv0;
    wire [31:0] c0_G16_mul0_G256_inv0;
    wire [31:0] c1_G16_mul0_G256_inv0;
    wire [31:0] d0_G16_mul0_G256_inv0;
    wire [31:0] d1_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G16_mul0_G256_inv0;
    wire [31:0] cxord_0_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G16_mul0_G256_inv0;
    wire [31:0] cxord_1_G16_mul0_G256_inv0;
    wire [31:0] r00_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r10_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3615_assgn3615;
    reg [31:0] z3615_assgn36150;
    reg [31:0] z3615_assgn36151;
    reg [31:0] z597_assgn597;
    wire [31:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3619_assgn3619;
    reg [31:0] z3619_assgn36190;
    reg [31:0] z3619_assgn36191;
    reg [31:0] z599_assgn599;
    wire [31:0] a1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3623_assgn3623;
    reg [31:0] z3623_assgn36230;
    reg [31:0] z3623_assgn36231;
    reg [31:0] z601_assgn601;
    wire [31:0] a0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3627_assgn3627;
    reg [31:0] z3627_assgn36270;
    reg [31:0] z3627_assgn36271;
    reg [31:0] z603_assgn603;
    wire [31:0] a1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3631_assgn3631;
    reg [31:0] z3631_assgn36310;
    reg [31:0] z3631_assgn36311;
    reg [31:0] z605_assgn605;
    wire [31:0] b0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3635_assgn3635;
    reg [31:0] z3635_assgn36350;
    reg [31:0] z3635_assgn36351;
    reg [31:0] z607_assgn607;
    wire [31:0] b1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] d0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] d1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] c0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] d0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] c1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] d1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] dec_2_inp_reg;
    wire [31:0] r0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3665_assgn3665;
    reg [31:0] z3665_assgn36650;
    reg [31:0] z635_assgn635;
    wire [31:0] u0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3669_assgn3669;
    reg [31:0] z3669_assgn36690;
    reg [31:0] z637_assgn637;
    wire [31:0] u1_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] cxord_0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] cxord_1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3677_assgn3677;
    reg [31:0] z3677_assgn36770;
    reg [31:0] z643_assgn643;
    wire [31:0] p0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] e0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3687_assgn3687;
    reg [31:0] z3687_assgn36870;
    reg [31:0] z651_assgn651;
    wire [31:0] p2_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] e1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3703_assgn3703;
    reg [31:0] z3703_assgn37030;
    reg [31:0] z665_assgn665;
    wire [31:0] u0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3707_assgn3707;
    reg [31:0] z3707_assgn37070;
    reg [31:0] z667_assgn667;
    wire [31:0] u1_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3711_assgn3711;
    reg [31:0] z3711_assgn37110;
    reg [31:0] z670_assgn670;
    reg [31:0] r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3715_assgn3715;
    reg [31:0] z3715_assgn37150;
    reg [31:0] z672_assgn672;
    wire [31:0] v1_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3719_assgn3719;
    reg [31:0] z3719_assgn37190;
    reg [31:0] z3719_assgn37191;
    reg [31:0] z673_assgn673;
    wire [31:0] p0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3729_assgn3729;
    reg [31:0] z3729_assgn37290;
    reg [31:0] z3729_assgn37291;
    reg [31:0] z681_assgn681;
    wire [31:0] p2_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3749_assgn3749;
    reg [31:0] z3749_assgn37490;
    reg [31:0] z699_assgn699;
    wire [31:0] u0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3753_assgn3753;
    reg [31:0] z3753_assgn37530;
    reg [31:0] z701_assgn701;
    wire [31:0] u1_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3757_assgn3757;
    reg [31:0] z3757_assgn37570;
    reg [31:0] z704_assgn704;
    reg [31:0] r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3761_assgn3761;
    reg [31:0] z3761_assgn37610;
    reg [31:0] z706_assgn706;
    wire [31:0] v1_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3765_assgn3765;
    reg [31:0] z3765_assgn37650;
    reg [31:0] z3765_assgn37651;
    reg [31:0] z707_assgn707;
    wire [31:0] p0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3775_assgn3775;
    reg [31:0] z3775_assgn37750;
    reg [31:0] z3775_assgn37751;
    reg [31:0] z715_assgn715;
    wire [31:0] p2_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3789_assgn3789;
    reg [31:0] z3789_assgn37890;
    reg [31:0] z3789_assgn37891;
    reg [31:0] z3789_assgn37892;
    reg [31:0] z727_assgn727;
    wire [31:0] p1ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z3793_assgn3793;
    reg [31:0] z3793_assgn37930;
    reg [31:0] z3793_assgn37931;
    reg [31:0] z3793_assgn37932;
    reg [31:0] z729_assgn729;
    wire [31:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] e0_G16_mul0_G256_inv0;
    wire [31:0] e1_G16_mul0_G256_inv0;
    wire [31:0] z3801_assgn3801;
    reg [31:0] z3801_assgn38010;
    reg [31:0] z3801_assgn38011;
    reg [31:0] z3801_assgn38012;
    reg [31:0] z735_assgn735;
    wire [31:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3805_assgn3805;
    reg [31:0] z3805_assgn38050;
    reg [31:0] z3805_assgn38051;
    reg [31:0] z3805_assgn38052;
    reg [31:0] z737_assgn737;
    wire [31:0] a1_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3809_assgn3809;
    reg [31:0] z3809_assgn38090;
    reg [31:0] z3809_assgn38091;
    reg [31:0] z3809_assgn38092;
    reg [31:0] z739_assgn739;
    wire [31:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3813_assgn3813;
    reg [31:0] z3813_assgn38130;
    reg [31:0] z3813_assgn38131;
    reg [31:0] z3813_assgn38132;
    reg [31:0] z741_assgn741;
    wire [31:0] a1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3817_assgn3817;
    reg [31:0] z3817_assgn38170;
    reg [31:0] z3817_assgn38171;
    reg [31:0] z3817_assgn38172;
    reg [31:0] z743_assgn743;
    wire [31:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3821_assgn3821;
    reg [31:0] z3821_assgn38210;
    reg [31:0] z3821_assgn38211;
    reg [31:0] z3821_assgn38212;
    reg [31:0] z745_assgn745;
    wire [31:0] b1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3833_assgn3833;
    reg [31:0] z3833_assgn38330;
    reg [31:0] z3833_assgn38331;
    reg [31:0] z3833_assgn38332;
    reg [31:0] z755_assgn755;
    wire [31:0] p1ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z3837_assgn3837;
    reg [31:0] z3837_assgn38370;
    reg [31:0] z3837_assgn38371;
    reg [31:0] z3837_assgn38372;
    reg [31:0] z757_assgn757;
    wire [31:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] e01_G16_mul0_G256_inv0;
    wire [31:0] e11_G16_mul0_G256_inv0;
    wire [31:0] r00_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r10_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3851_assgn3851;
    reg [31:0] z3851_assgn38510;
    reg [31:0] z3851_assgn38511;
    reg [31:0] z769_assgn769;
    wire [31:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3855_assgn3855;
    reg [31:0] z3855_assgn38550;
    reg [31:0] z3855_assgn38551;
    reg [31:0] z771_assgn771;
    wire [31:0] a1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3859_assgn3859;
    reg [31:0] z3859_assgn38590;
    reg [31:0] z3859_assgn38591;
    reg [31:0] z773_assgn773;
    wire [31:0] a0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3863_assgn3863;
    reg [31:0] z3863_assgn38630;
    reg [31:0] z3863_assgn38631;
    reg [31:0] z775_assgn775;
    wire [31:0] a1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3867_assgn3867;
    reg [31:0] z3867_assgn38670;
    reg [31:0] z3867_assgn38671;
    reg [31:0] z777_assgn777;
    wire [31:0] b0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3871_assgn3871;
    reg [31:0] z3871_assgn38710;
    reg [31:0] z3871_assgn38711;
    reg [31:0] z779_assgn779;
    wire [31:0] b1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] d0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] d1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] c0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] d0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] c1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] d1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3901_assgn3901;
    reg [31:0] z3901_assgn39010;
    reg [31:0] z807_assgn807;
    wire [31:0] u0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3905_assgn3905;
    reg [31:0] z3905_assgn39050;
    reg [31:0] z809_assgn809;
    wire [31:0] u1_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] cxord_0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] cxord_1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3913_assgn3913;
    reg [31:0] z3913_assgn39130;
    reg [31:0] z815_assgn815;
    wire [31:0] p0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] e0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3923_assgn3923;
    reg [31:0] z3923_assgn39230;
    reg [31:0] z823_assgn823;
    wire [31:0] p2_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] e1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3939_assgn3939;
    reg [31:0] z3939_assgn39390;
    reg [31:0] z837_assgn837;
    wire [31:0] u0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3943_assgn3943;
    reg [31:0] z3943_assgn39430;
    reg [31:0] z839_assgn839;
    wire [31:0] u1_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3947_assgn3947;
    reg [31:0] z3947_assgn39470;
    reg [31:0] z842_assgn842;
    reg [31:0] r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3951_assgn3951;
    reg [31:0] z3951_assgn39510;
    reg [31:0] z844_assgn844;
    wire [31:0] v1_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3955_assgn3955;
    reg [31:0] z3955_assgn39550;
    reg [31:0] z3955_assgn39551;
    reg [31:0] z845_assgn845;
    wire [31:0] p0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3965_assgn3965;
    reg [31:0] z3965_assgn39650;
    reg [31:0] z3965_assgn39651;
    reg [31:0] z853_assgn853;
    wire [31:0] p2_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3985_assgn3985;
    reg [31:0] z3985_assgn39850;
    reg [31:0] z871_assgn871;
    wire [31:0] u0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3989_assgn3989;
    reg [31:0] z3989_assgn39890;
    reg [31:0] z873_assgn873;
    wire [31:0] u1_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3993_assgn3993;
    reg [31:0] z3993_assgn39930;
    reg [31:0] z876_assgn876;
    reg [31:0] r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z3997_assgn3997;
    reg [31:0] z3997_assgn39970;
    reg [31:0] z878_assgn878;
    wire [31:0] v1_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z4001_assgn4001;
    reg [31:0] z4001_assgn40010;
    reg [31:0] z4001_assgn40011;
    reg [31:0] z879_assgn879;
    wire [31:0] p0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z4011_assgn4011;
    reg [31:0] z4011_assgn40110;
    reg [31:0] z4011_assgn40111;
    reg [31:0] z887_assgn887;
    wire [31:0] p2_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z4025_assgn4025;
    reg [31:0] z4025_assgn40250;
    reg [31:0] z4025_assgn40251;
    reg [31:0] z4025_assgn40252;
    reg [31:0] z899_assgn899;
    wire [31:0] p1ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z4029_assgn4029;
    reg [31:0] z4029_assgn40290;
    reg [31:0] z4029_assgn40291;
    reg [31:0] z4029_assgn40292;
    reg [31:0] z901_assgn901;
    wire [31:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p0_0_G16_mul0_G256_inv0;
    wire [31:0] p1_0_G16_mul0_G256_inv0;
    wire [31:0] p0_G16_mul0_G256_inv0;
    wire [31:0] p1_G16_mul0_G256_inv0;
    wire [31:0] r00_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r10_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4047_assgn4047;
    reg [31:0] z4047_assgn40470;
    reg [31:0] z4047_assgn40471;
    reg [31:0] z917_assgn917;
    wire [31:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4051_assgn4051;
    reg [31:0] z4051_assgn40510;
    reg [31:0] z4051_assgn40511;
    reg [31:0] z919_assgn919;
    wire [31:0] a1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4055_assgn4055;
    reg [31:0] z4055_assgn40550;
    reg [31:0] z4055_assgn40551;
    reg [31:0] z921_assgn921;
    wire [31:0] a0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4059_assgn4059;
    reg [31:0] z4059_assgn40590;
    reg [31:0] z4059_assgn40591;
    reg [31:0] z923_assgn923;
    wire [31:0] a1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4063_assgn4063;
    reg [31:0] z4063_assgn40630;
    reg [31:0] z4063_assgn40631;
    reg [31:0] z925_assgn925;
    wire [31:0] b0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4067_assgn4067;
    reg [31:0] z4067_assgn40670;
    reg [31:0] z4067_assgn40671;
    reg [31:0] z927_assgn927;
    wire [31:0] b1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] d0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] d1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] c0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] d0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] c1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] d1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4097_assgn4097;
    reg [31:0] z4097_assgn40970;
    reg [31:0] z955_assgn955;
    wire [31:0] u0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4101_assgn4101;
    reg [31:0] z4101_assgn41010;
    reg [31:0] z957_assgn957;
    wire [31:0] u1_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] cxord_0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] cxord_1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4109_assgn4109;
    reg [31:0] z4109_assgn41090;
    reg [31:0] z963_assgn963;
    wire [31:0] p0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] e0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4119_assgn4119;
    reg [31:0] z4119_assgn41190;
    reg [31:0] z971_assgn971;
    wire [31:0] p2_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] e1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4135_assgn4135;
    reg [31:0] z4135_assgn41350;
    reg [31:0] z985_assgn985;
    wire [31:0] u0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4139_assgn4139;
    reg [31:0] z4139_assgn41390;
    reg [31:0] z987_assgn987;
    wire [31:0] u1_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4143_assgn4143;
    reg [31:0] z4143_assgn41430;
    reg [31:0] z990_assgn990;
    reg [31:0] r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4147_assgn4147;
    reg [31:0] z4147_assgn41470;
    reg [31:0] z992_assgn992;
    wire [31:0] v1_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4151_assgn4151;
    reg [31:0] z4151_assgn41510;
    reg [31:0] z4151_assgn41511;
    reg [31:0] z993_assgn993;
    wire [31:0] p0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4161_assgn4161;
    reg [31:0] z4161_assgn41610;
    reg [31:0] z4161_assgn41611;
    reg [31:0] z1001_assgn1001;
    wire [31:0] p2_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4181_assgn4181;
    reg [31:0] z4181_assgn41810;
    reg [31:0] z1019_assgn1019;
    wire [31:0] u0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4185_assgn4185;
    reg [31:0] z4185_assgn41850;
    reg [31:0] z1021_assgn1021;
    wire [31:0] u1_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4189_assgn4189;
    reg [31:0] z4189_assgn41890;
    reg [31:0] z1024_assgn1024;
    reg [31:0] r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4193_assgn4193;
    reg [31:0] z4193_assgn41930;
    reg [31:0] z1026_assgn1026;
    wire [31:0] v1_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4197_assgn4197;
    reg [31:0] z4197_assgn41970;
    reg [31:0] z4197_assgn41971;
    reg [31:0] z1027_assgn1027;
    wire [31:0] p0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4207_assgn4207;
    reg [31:0] z4207_assgn42070;
    reg [31:0] z4207_assgn42071;
    reg [31:0] z1035_assgn1035;
    wire [31:0] p2_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4221_assgn4221;
    reg [31:0] z4221_assgn42210;
    reg [31:0] z4221_assgn42211;
    reg [31:0] z4221_assgn42212;
    reg [31:0] z1047_assgn1047;
    wire [31:0] p1ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4225_assgn4225;
    reg [31:0] z4225_assgn42250;
    reg [31:0] z4225_assgn42251;
    reg [31:0] z4225_assgn42252;
    reg [31:0] z1049_assgn1049;
    wire [31:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q0_0_G16_mul0_G256_inv0;
    wire [31:0] q1_0_G16_mul0_G256_inv0;
    wire [31:0] q0_G16_mul0_G256_inv0;
    wire [31:0] q1_G16_mul0_G256_inv0;
    wire [31:0] z4237_assgn4237;
    reg [31:0] z4237_assgn42370;
    reg [31:0] z4237_assgn42371;
    reg [31:0] z4237_assgn42372;
    reg [31:0] z1059_assgn1059;
    wire [31:0] p0ls2_G16_mul0_G256_inv0;
    wire [31:0] z4241_assgn4241;
    reg [31:0] z4241_assgn42410;
    reg [31:0] z4241_assgn42411;
    reg [31:0] z4241_assgn42412;
    reg [31:0] z1061_assgn1061;
    wire [31:0] p1ls2_G16_mul0_G256_inv0;
    wire [31:0] d0_G256_inv0;
    wire [31:0] d1_G256_inv0;
    wire [31:0] c0xord0_G256_inv0;
    wire [31:0] c1xord1_G256_inv0;
    wire [31:0] z4253_assgn4253;
    reg [31:0] z4253_assgn42530;
    reg [31:0] z4253_assgn42531;
    reg [31:0] z4253_assgn42532;
    reg [31:0] z1071_assgn1071;
    wire [31:0] r00_G16_inv0_G256_inv0;
    wire [31:0] z4257_assgn4257;
    reg [31:0] z4257_assgn42570;
    reg [31:0] z4257_assgn42571;
    reg [31:0] z4257_assgn42572;
    reg [31:0] z1073_assgn1073;
    wire [31:0] r10_G16_inv0_G256_inv0;
    wire [31:0] z4261_assgn4261;
    reg [31:0] z4261_assgn42610;
    reg [31:0] z4261_assgn42611;
    reg [31:0] z4261_assgn42612;
    reg [31:0] z1075_assgn1075;
    wire [31:0] r20_G16_inv0_G256_inv0;
    wire [31:0] z4265_assgn4265;
    reg [31:0] z4265_assgn42650;
    reg [31:0] z4265_assgn42651;
    reg [31:0] z4265_assgn42652;
    reg [31:0] z4265_assgn42653;
    reg [31:0] z1077_assgn1077;
    wire [31:0] r30_G16_inv0_G256_inv0;
    wire [31:0] z4269_assgn4269;
    reg [31:0] z4269_assgn42690;
    reg [31:0] z4269_assgn42691;
    reg [31:0] z4269_assgn42692;
    reg [31:0] z4269_assgn42693;
    reg [31:0] z1079_assgn1079;
    wire [31:0] r40_G16_inv0_G256_inv0;
    wire [31:0] z4273_assgn4273;
    reg [31:0] z4273_assgn42730;
    reg [31:0] z4273_assgn42731;
    reg [31:0] z4273_assgn42732;
    reg [31:0] z4273_assgn42733;
    reg [31:0] z1081_assgn1081;
    wire [31:0] r50_G16_inv0_G256_inv0;
    wire [31:0] z4277_assgn4277;
    reg [31:0] z4277_assgn42770;
    reg [31:0] z4277_assgn42771;
    reg [31:0] z4277_assgn42772;
    reg [31:0] z4277_assgn42773;
    reg [31:0] z1083_assgn1083;
    wire [31:0] r60_G16_inv0_G256_inv0;
    wire [31:0] z4281_assgn4281;
    reg [31:0] z4281_assgn42810;
    reg [31:0] z4281_assgn42811;
    reg [31:0] z4281_assgn42812;
    reg [31:0] z4281_assgn42813;
    reg [31:0] z1085_assgn1085;
    wire [31:0] r70_G16_inv0_G256_inv0;
    wire [31:0] z4285_assgn4285;
    reg [31:0] z4285_assgn42850;
    reg [31:0] z4285_assgn42851;
    reg [31:0] z4285_assgn42852;
    reg [31:0] z4285_assgn42853;
    reg [31:0] z1087_assgn1087;
    wire [31:0] r80_G16_inv0_G256_inv0;
    wire [31:0] z4289_assgn4289;
    reg [31:0] z4289_assgn42890;
    reg [31:0] z4289_assgn42891;
    reg [31:0] z4289_assgn42892;
    reg [31:0] z4289_assgn42893;
    reg [31:0] z1089_assgn1089;
    reg [31:0] c0xord0_G256_inv0_reg;
    wire [31:0] a0_0_G16_inv0_G256_inv0;
    wire [31:0] z4293_assgn4293;
    reg [31:0] z4293_assgn42930;
    reg [31:0] z4293_assgn42931;
    reg [31:0] z4293_assgn42932;
    reg [31:0] z4293_assgn42933;
    reg [31:0] z1091_assgn1091;
    reg [31:0] c1xord1_G256_inv0_reg;
    wire [31:0] a1_0_G16_inv0_G256_inv0;
    wire [31:0] z4297_assgn4297;
    reg [31:0] z4297_assgn42970;
    reg [31:0] z4297_assgn42971;
    reg [31:0] z4297_assgn42972;
    reg [31:0] z4297_assgn42973;
    reg [31:0] z1093_assgn1093;
    wire [31:0] a0_G16_inv0_G256_inv0;
    wire [31:0] z4301_assgn4301;
    reg [31:0] z4301_assgn43010;
    reg [31:0] z4301_assgn43011;
    reg [31:0] z4301_assgn43012;
    reg [31:0] z4301_assgn43013;
    reg [31:0] z1095_assgn1095;
    wire [31:0] a1_G16_inv0_G256_inv0;
    wire [31:0] z4305_assgn4305;
    reg [31:0] z4305_assgn43050;
    reg [31:0] z4305_assgn43051;
    reg [31:0] z4305_assgn43052;
    reg [31:0] z1097_assgn1097;
    wire [31:0] b0_G16_inv0_G256_inv0;
    wire [31:0] z4309_assgn4309;
    reg [31:0] z4309_assgn43090;
    reg [31:0] z4309_assgn43091;
    reg [31:0] z4309_assgn43092;
    reg [31:0] z1099_assgn1099;
    wire [31:0] b1_G16_inv0_G256_inv0;
    wire [31:0] z4313_assgn4313;
    reg [31:0] z4313_assgn43130;
    reg [31:0] z4313_assgn43131;
    reg [31:0] z4313_assgn43132;
    reg [31:0] z1101_assgn1101;
    wire [31:0] z4315_assgn4315;
    reg [31:0] z4315_assgn43150;
    reg [31:0] z4315_assgn43151;
    reg [31:0] z1102_assgn1102;
    wire [31:0] a0xorb0_G16_inv0_G256_inv0;
    wire [31:0] z4319_assgn4319;
    reg [31:0] z4319_assgn43190;
    reg [31:0] z4319_assgn43191;
    reg [31:0] z4319_assgn43192;
    reg [31:0] z1103_assgn1103;
    wire [31:0] z4321_assgn4321;
    reg [31:0] z4321_assgn43210;
    reg [31:0] z4321_assgn43211;
    reg [31:0] z1104_assgn1104;
    wire [31:0] a1xorb1_G16_inv0_G256_inv0;
    wire [31:0] z4325_assgn4325;
    reg [31:0] z4325_assgn43250;
    reg [31:0] z4325_assgn43251;
    reg [31:0] z4325_assgn43252;
    reg [31:0] z4325_assgn43253;
    reg [31:0] z4325_assgn43254;
    reg [31:0] z4325_assgn43255;
    reg [31:0] z4325_assgn43256;
    reg [31:0] z1105_assgn1105;
    wire [31:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4329_assgn4329;
    reg [31:0] z4329_assgn43290;
    reg [31:0] z4329_assgn43291;
    reg [31:0] z4329_assgn43292;
    reg [31:0] z4329_assgn43293;
    reg [31:0] z4329_assgn43294;
    reg [31:0] z4329_assgn43295;
    reg [31:0] z4329_assgn43296;
    reg [31:0] z1107_assgn1107;
    wire [31:0] a1_0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4333_assgn4333;
    reg [31:0] z4333_assgn43330;
    reg [31:0] z4333_assgn43331;
    reg [31:0] z4333_assgn43332;
    reg [31:0] z4333_assgn43333;
    reg [31:0] z4333_assgn43334;
    reg [31:0] z4333_assgn43335;
    reg [31:0] z4333_assgn43336;
    reg [31:0] z1109_assgn1109;
    wire [31:0] a0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4337_assgn4337;
    reg [31:0] z4337_assgn43370;
    reg [31:0] z4337_assgn43371;
    reg [31:0] z4337_assgn43372;
    reg [31:0] z4337_assgn43373;
    reg [31:0] z4337_assgn43374;
    reg [31:0] z4337_assgn43375;
    reg [31:0] z4337_assgn43376;
    reg [31:0] z1111_assgn1111;
    wire [31:0] a1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4341_assgn4341;
    reg [31:0] z4341_assgn43410;
    reg [31:0] z4341_assgn43411;
    reg [31:0] z4341_assgn43412;
    reg [31:0] z4341_assgn43413;
    reg [31:0] z4341_assgn43414;
    reg [31:0] z4341_assgn43415;
    reg [31:0] z4341_assgn43416;
    reg [31:0] z1113_assgn1113;
    wire [31:0] b0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4345_assgn4345;
    reg [31:0] z4345_assgn43450;
    reg [31:0] z4345_assgn43451;
    reg [31:0] z4345_assgn43452;
    reg [31:0] z4345_assgn43453;
    reg [31:0] z4345_assgn43454;
    reg [31:0] z4345_assgn43455;
    reg [31:0] z4345_assgn43456;
    reg [31:0] z1115_assgn1115;
    wire [31:0] b1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4349_assgn4349;
    reg [31:0] z4349_assgn43490;
    reg [31:0] z4349_assgn43491;
    reg [31:0] z4349_assgn43492;
    reg [31:0] z4349_assgn43493;
    reg [31:0] z4349_assgn43494;
    reg [31:0] z4349_assgn43495;
    reg [31:0] z4349_assgn43496;
    reg [31:0] z1117_assgn1117;
    wire [31:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4353_assgn4353;
    reg [31:0] z4353_assgn43530;
    reg [31:0] z4353_assgn43531;
    reg [31:0] z4353_assgn43532;
    reg [31:0] z4353_assgn43533;
    reg [31:0] z4353_assgn43534;
    reg [31:0] z4353_assgn43535;
    reg [31:0] z4353_assgn43536;
    reg [31:0] z1119_assgn1119;
    wire [31:0] b1ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] c0_0_G16_inv0_G256_inv0;
    wire [31:0] c1_0_G16_inv0_G256_inv0;
    wire [31:0] z4361_assgn4361;
    reg [31:0] z4361_assgn43610;
    reg [31:0] z4361_assgn43611;
    reg [31:0] z4361_assgn43612;
    reg [31:0] z4361_assgn43613;
    reg [31:0] z4361_assgn43614;
    reg [31:0] z4361_assgn43615;
    reg [31:0] z4361_assgn43616;
    reg [31:0] z1125_assgn1125;
    wire [31:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4365_assgn4365;
    reg [31:0] z4365_assgn43650;
    reg [31:0] z4365_assgn43651;
    reg [31:0] z4365_assgn43652;
    reg [31:0] z4365_assgn43653;
    reg [31:0] z4365_assgn43654;
    reg [31:0] z4365_assgn43655;
    reg [31:0] z4365_assgn43656;
    reg [31:0] z1127_assgn1127;
    wire [31:0] a1_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4369_assgn4369;
    reg [31:0] z4369_assgn43690;
    reg [31:0] z4369_assgn43691;
    reg [31:0] z4369_assgn43692;
    reg [31:0] z4369_assgn43693;
    reg [31:0] z4369_assgn43694;
    reg [31:0] z4369_assgn43695;
    reg [31:0] z4369_assgn43696;
    reg [31:0] z1129_assgn1129;
    wire [31:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4373_assgn4373;
    reg [31:0] z4373_assgn43730;
    reg [31:0] z4373_assgn43731;
    reg [31:0] z4373_assgn43732;
    reg [31:0] z4373_assgn43733;
    reg [31:0] z4373_assgn43734;
    reg [31:0] z4373_assgn43735;
    reg [31:0] z4373_assgn43736;
    reg [31:0] z1131_assgn1131;
    wire [31:0] a1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4377_assgn4377;
    reg [31:0] z4377_assgn43770;
    reg [31:0] z4377_assgn43771;
    reg [31:0] z4377_assgn43772;
    reg [31:0] z4377_assgn43773;
    reg [31:0] z4377_assgn43774;
    reg [31:0] z4377_assgn43775;
    reg [31:0] z4377_assgn43776;
    reg [31:0] z1133_assgn1133;
    wire [31:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4381_assgn4381;
    reg [31:0] z4381_assgn43810;
    reg [31:0] z4381_assgn43811;
    reg [31:0] z4381_assgn43812;
    reg [31:0] z4381_assgn43813;
    reg [31:0] z4381_assgn43814;
    reg [31:0] z4381_assgn43815;
    reg [31:0] z4381_assgn43816;
    reg [31:0] z1135_assgn1135;
    wire [31:0] b1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4393_assgn4393;
    reg [31:0] z4393_assgn43930;
    reg [31:0] z4393_assgn43931;
    reg [31:0] z4393_assgn43932;
    reg [31:0] z4393_assgn43933;
    reg [31:0] z4393_assgn43934;
    reg [31:0] z4393_assgn43935;
    reg [31:0] z4393_assgn43936;
    reg [31:0] z1145_assgn1145;
    wire [31:0] p1ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4397_assgn4397;
    reg [31:0] z4397_assgn43970;
    reg [31:0] z4397_assgn43971;
    reg [31:0] z4397_assgn43972;
    reg [31:0] z4397_assgn43973;
    reg [31:0] z4397_assgn43974;
    reg [31:0] z4397_assgn43975;
    reg [31:0] z4397_assgn43976;
    reg [31:0] z1147_assgn1147;
    wire [31:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] c0_G16_inv0_G256_inv0;
    wire [31:0] c1_G16_inv0_G256_inv0;
    wire [31:0] z4405_assgn4405;
    reg [31:0] z4405_assgn44050;
    reg [31:0] z4405_assgn44051;
    reg [31:0] z4405_assgn44052;
    reg [31:0] z1153_assgn1153;
    wire [31:0] r00_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4409_assgn4409;
    reg [31:0] z4409_assgn44090;
    reg [31:0] z4409_assgn44091;
    reg [31:0] z4409_assgn44092;
    reg [31:0] z1155_assgn1155;
    wire [31:0] r10_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4413_assgn4413;
    reg [31:0] z4413_assgn44130;
    reg [31:0] z4413_assgn44131;
    reg [31:0] z4413_assgn44132;
    reg [31:0] z1157_assgn1157;
    wire [31:0] r20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4417_assgn4417;
    reg [31:0] z4417_assgn44170;
    reg [31:0] z4417_assgn44171;
    reg [31:0] z4417_assgn44172;
    reg [31:0] z4417_assgn44173;
    reg [31:0] z4417_assgn44174;
    reg [31:0] z4417_assgn44175;
    reg [31:0] z1159_assgn1159;
    wire [31:0] z4419_assgn4419;
    reg [31:0] z4419_assgn44190;
    reg [31:0] z1160_assgn1160;
    wire [31:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4423_assgn4423;
    reg [31:0] z4423_assgn44230;
    reg [31:0] z4423_assgn44231;
    reg [31:0] z4423_assgn44232;
    reg [31:0] z4423_assgn44233;
    reg [31:0] z4423_assgn44234;
    reg [31:0] z4423_assgn44235;
    reg [31:0] z1161_assgn1161;
    wire [31:0] z4425_assgn4425;
    reg [31:0] z4425_assgn44250;
    reg [31:0] z1162_assgn1162;
    wire [31:0] a1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4429_assgn4429;
    reg [31:0] z4429_assgn44290;
    reg [31:0] z4429_assgn44291;
    reg [31:0] z4429_assgn44292;
    reg [31:0] z4429_assgn44293;
    reg [31:0] z4429_assgn44294;
    reg [31:0] z4429_assgn44295;
    reg [31:0] z1163_assgn1163;
    wire [31:0] a0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4433_assgn4433;
    reg [31:0] z4433_assgn44330;
    reg [31:0] z4433_assgn44331;
    reg [31:0] z4433_assgn44332;
    reg [31:0] z4433_assgn44333;
    reg [31:0] z4433_assgn44334;
    reg [31:0] z4433_assgn44335;
    reg [31:0] z1165_assgn1165;
    wire [31:0] a1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4437_assgn4437;
    reg [31:0] z4437_assgn44370;
    reg [31:0] z4437_assgn44371;
    reg [31:0] z4437_assgn44372;
    reg [31:0] z4437_assgn44373;
    reg [31:0] z4437_assgn44374;
    reg [31:0] z4437_assgn44375;
    reg [31:0] z1167_assgn1167;
    wire [31:0] z4439_assgn4439;
    reg [31:0] z4439_assgn44390;
    reg [31:0] z1168_assgn1168;
    wire [31:0] b0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4443_assgn4443;
    reg [31:0] z4443_assgn44430;
    reg [31:0] z4443_assgn44431;
    reg [31:0] z4443_assgn44432;
    reg [31:0] z4443_assgn44433;
    reg [31:0] z4443_assgn44434;
    reg [31:0] z4443_assgn44435;
    reg [31:0] z1169_assgn1169;
    wire [31:0] z4445_assgn4445;
    reg [31:0] z4445_assgn44450;
    reg [31:0] z1170_assgn1170;
    wire [31:0] b1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4449_assgn4449;
    reg [31:0] z4449_assgn44490;
    reg [31:0] z4449_assgn44491;
    reg [31:0] z4449_assgn44492;
    reg [31:0] z1171_assgn1171;
    wire [31:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4453_assgn4453;
    reg [31:0] z4453_assgn44530;
    reg [31:0] z4453_assgn44531;
    reg [31:0] z4453_assgn44532;
    reg [31:0] z1173_assgn1173;
    wire [31:0] c1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4457_assgn4457;
    reg [31:0] z4457_assgn44570;
    reg [31:0] z4457_assgn44571;
    reg [31:0] z4457_assgn44572;
    reg [31:0] z1175_assgn1175;
    wire [31:0] c0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4461_assgn4461;
    reg [31:0] z4461_assgn44610;
    reg [31:0] z4461_assgn44611;
    reg [31:0] z4461_assgn44612;
    reg [31:0] z1177_assgn1177;
    wire [31:0] c1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4465_assgn4465;
    reg [31:0] z4465_assgn44650;
    reg [31:0] z4465_assgn44651;
    reg [31:0] z4465_assgn44652;
    reg [31:0] z1179_assgn1179;
    wire [31:0] d0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4469_assgn4469;
    reg [31:0] z4469_assgn44690;
    reg [31:0] z4469_assgn44691;
    reg [31:0] z4469_assgn44692;
    reg [31:0] z1181_assgn1181;
    wire [31:0] d1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] c0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] d0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] axorb_1_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] c1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] d1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4481_assgn4481;
    reg [31:0] z4481_assgn44810;
    reg [31:0] z4481_assgn44811;
    reg [31:0] z4481_assgn44812;
    reg [31:0] z4481_assgn44813;
    reg [31:0] z1191_assgn1191;
    wire [31:0] r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4489_assgn4489;
    reg [31:0] z4489_assgn44890;
    reg [31:0] z1197_assgn1197;
    wire [31:0] u0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4493_assgn4493;
    reg [31:0] z4493_assgn44930;
    reg [31:0] z1199_assgn1199;
    wire [31:0] u1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] cxord_0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] cxord_1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4501_assgn4501;
    reg [31:0] z4501_assgn45010;
    reg [31:0] z1205_assgn1205;
    wire [31:0] p0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] e0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4511_assgn4511;
    reg [31:0] z4511_assgn45110;
    reg [31:0] z1213_assgn1213;
    wire [31:0] p2_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] e1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4521_assgn4521;
    reg [31:0] z4521_assgn45210;
    reg [31:0] z4521_assgn45211;
    reg [31:0] z4521_assgn45212;
    reg [31:0] z4521_assgn45213;
    reg [31:0] z1221_assgn1221;
    wire [31:0] r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4529_assgn4529;
    reg [31:0] z4529_assgn45290;
    reg [31:0] z1227_assgn1227;
    wire [31:0] u0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4533_assgn4533;
    reg [31:0] z4533_assgn45330;
    reg [31:0] z1229_assgn1229;
    wire [31:0] u1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4537_assgn4537;
    reg [31:0] z4537_assgn45370;
    reg [31:0] z1232_assgn1232;
    reg [31:0] r0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4541_assgn4541;
    reg [31:0] z4541_assgn45410;
    reg [31:0] z1234_assgn1234;
    wire [31:0] v1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4545_assgn4545;
    reg [31:0] z4545_assgn45450;
    reg [31:0] z4545_assgn45451;
    reg [31:0] z1235_assgn1235;
    wire [31:0] p0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4555_assgn4555;
    reg [31:0] z4555_assgn45550;
    reg [31:0] z4555_assgn45551;
    reg [31:0] z1243_assgn1243;
    wire [31:0] p2_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4569_assgn4569;
    reg [31:0] z4569_assgn45690;
    reg [31:0] z4569_assgn45691;
    reg [31:0] z4569_assgn45692;
    reg [31:0] z4569_assgn45693;
    reg [31:0] z1255_assgn1255;
    wire [31:0] r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4577_assgn4577;
    reg [31:0] z4577_assgn45770;
    reg [31:0] z1261_assgn1261;
    wire [31:0] u0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4581_assgn4581;
    reg [31:0] z4581_assgn45810;
    reg [31:0] z1263_assgn1263;
    wire [31:0] u1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4585_assgn4585;
    reg [31:0] z4585_assgn45850;
    reg [31:0] z1266_assgn1266;
    reg [31:0] r0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4589_assgn4589;
    reg [31:0] z4589_assgn45890;
    reg [31:0] z1268_assgn1268;
    wire [31:0] v1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4593_assgn4593;
    reg [31:0] z4593_assgn45930;
    reg [31:0] z4593_assgn45931;
    reg [31:0] z1269_assgn1269;
    wire [31:0] p0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4603_assgn4603;
    reg [31:0] z4603_assgn46030;
    reg [31:0] z4603_assgn46031;
    reg [31:0] z1277_assgn1277;
    wire [31:0] p2_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4617_assgn4617;
    reg [31:0] z4617_assgn46170;
    reg [31:0] z4617_assgn46171;
    reg [31:0] z4617_assgn46172;
    reg [31:0] z4617_assgn46173;
    reg [31:0] z4617_assgn46174;
    reg [31:0] z4617_assgn46175;
    reg [31:0] z4617_assgn46176;
    reg [31:0] z1289_assgn1289;
    wire [31:0] p1ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4621_assgn4621;
    reg [31:0] z4621_assgn46210;
    reg [31:0] z4621_assgn46211;
    reg [31:0] z4621_assgn46212;
    reg [31:0] z4621_assgn46213;
    reg [31:0] z4621_assgn46214;
    reg [31:0] z4621_assgn46215;
    reg [31:0] z4621_assgn46216;
    reg [31:0] z1291_assgn1291;
    wire [31:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] d0_G16_inv0_G256_inv0;
    wire [31:0] d1_G16_inv0_G256_inv0;
    wire [31:0] c0xord0_G16_inv0_G256_inv0;
    wire [31:0] c1xord1_G16_inv0_G256_inv0;
    wire [31:0] z4633_assgn4633;
    reg [31:0] z4633_assgn46330;
    reg [31:0] z4633_assgn46331;
    reg [31:0] z4633_assgn46332;
    reg [31:0] z4633_assgn46333;
    reg [31:0] z4633_assgn46334;
    reg [31:0] z4633_assgn46335;
    reg [31:0] z4633_assgn46336;
    reg [31:0] z1301_assgn1301;
    wire [31:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4637_assgn4637;
    reg [31:0] z4637_assgn46370;
    reg [31:0] z4637_assgn46371;
    reg [31:0] z4637_assgn46372;
    reg [31:0] z4637_assgn46373;
    reg [31:0] z4637_assgn46374;
    reg [31:0] z4637_assgn46375;
    reg [31:0] z4637_assgn46376;
    reg [31:0] z1303_assgn1303;
    wire [31:0] a1_0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4641_assgn4641;
    reg [31:0] z4641_assgn46410;
    reg [31:0] z4641_assgn46411;
    reg [31:0] z4641_assgn46412;
    reg [31:0] z4641_assgn46413;
    reg [31:0] z4641_assgn46414;
    reg [31:0] z4641_assgn46415;
    reg [31:0] z4641_assgn46416;
    reg [31:0] z1305_assgn1305;
    wire [31:0] a0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4645_assgn4645;
    reg [31:0] z4645_assgn46450;
    reg [31:0] z4645_assgn46451;
    reg [31:0] z4645_assgn46452;
    reg [31:0] z4645_assgn46453;
    reg [31:0] z4645_assgn46454;
    reg [31:0] z4645_assgn46455;
    reg [31:0] z4645_assgn46456;
    reg [31:0] z1307_assgn1307;
    wire [31:0] a1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4649_assgn4649;
    reg [31:0] z4649_assgn46490;
    reg [31:0] z4649_assgn46491;
    reg [31:0] z4649_assgn46492;
    reg [31:0] z4649_assgn46493;
    reg [31:0] z4649_assgn46494;
    reg [31:0] z4649_assgn46495;
    reg [31:0] z4649_assgn46496;
    reg [31:0] z1309_assgn1309;
    wire [31:0] b0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4653_assgn4653;
    reg [31:0] z4653_assgn46530;
    reg [31:0] z4653_assgn46531;
    reg [31:0] z4653_assgn46532;
    reg [31:0] z4653_assgn46533;
    reg [31:0] z4653_assgn46534;
    reg [31:0] z4653_assgn46535;
    reg [31:0] z4653_assgn46536;
    reg [31:0] z1311_assgn1311;
    wire [31:0] b1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4657_assgn4657;
    reg [31:0] z4657_assgn46570;
    reg [31:0] z4657_assgn46571;
    reg [31:0] z4657_assgn46572;
    reg [31:0] z4657_assgn46573;
    reg [31:0] z4657_assgn46574;
    reg [31:0] z4657_assgn46575;
    reg [31:0] z4657_assgn46576;
    reg [31:0] z1313_assgn1313;
    wire [31:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z4661_assgn4661;
    reg [31:0] z4661_assgn46610;
    reg [31:0] z4661_assgn46611;
    reg [31:0] z4661_assgn46612;
    reg [31:0] z4661_assgn46613;
    reg [31:0] z4661_assgn46614;
    reg [31:0] z4661_assgn46615;
    reg [31:0] z4661_assgn46616;
    reg [31:0] z1315_assgn1315;
    wire [31:0] b1ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] e0_G16_inv0_G256_inv0;
    wire [31:0] e1_G16_inv0_G256_inv0;
    wire [31:0] z4669_assgn4669;
    reg [31:0] z4669_assgn46690;
    reg [31:0] z4669_assgn46691;
    reg [31:0] z4669_assgn46692;
    reg [31:0] z4669_assgn46693;
    reg [31:0] z1321_assgn1321;
    wire [31:0] r00_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4673_assgn4673;
    reg [31:0] z4673_assgn46730;
    reg [31:0] z4673_assgn46731;
    reg [31:0] z4673_assgn46732;
    reg [31:0] z4673_assgn46733;
    reg [31:0] z1323_assgn1323;
    wire [31:0] r10_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4677_assgn4677;
    reg [31:0] z4677_assgn46770;
    reg [31:0] z4677_assgn46771;
    reg [31:0] z4677_assgn46772;
    reg [31:0] z4677_assgn46773;
    reg [31:0] z1325_assgn1325;
    wire [31:0] r20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4681_assgn4681;
    reg [31:0] z4681_assgn46810;
    reg [31:0] z4681_assgn46811;
    reg [31:0] z4681_assgn46812;
    reg [31:0] z4681_assgn46813;
    reg [31:0] z4681_assgn46814;
    reg [31:0] z4681_assgn46815;
    reg [31:0] z4681_assgn46816;
    reg [31:0] z1327_assgn1327;
    wire [31:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4685_assgn4685;
    reg [31:0] z4685_assgn46850;
    reg [31:0] z4685_assgn46851;
    reg [31:0] z4685_assgn46852;
    reg [31:0] z4685_assgn46853;
    reg [31:0] z4685_assgn46854;
    reg [31:0] z4685_assgn46855;
    reg [31:0] z4685_assgn46856;
    reg [31:0] z1329_assgn1329;
    wire [31:0] a1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4689_assgn4689;
    reg [31:0] z4689_assgn46890;
    reg [31:0] z4689_assgn46891;
    reg [31:0] z4689_assgn46892;
    reg [31:0] z4689_assgn46893;
    reg [31:0] z4689_assgn46894;
    reg [31:0] z4689_assgn46895;
    reg [31:0] z4689_assgn46896;
    reg [31:0] z1331_assgn1331;
    wire [31:0] a0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4693_assgn4693;
    reg [31:0] z4693_assgn46930;
    reg [31:0] z4693_assgn46931;
    reg [31:0] z4693_assgn46932;
    reg [31:0] z4693_assgn46933;
    reg [31:0] z4693_assgn46934;
    reg [31:0] z4693_assgn46935;
    reg [31:0] z4693_assgn46936;
    reg [31:0] z1333_assgn1333;
    wire [31:0] a1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4697_assgn4697;
    reg [31:0] z4697_assgn46970;
    reg [31:0] z4697_assgn46971;
    reg [31:0] z4697_assgn46972;
    reg [31:0] z4697_assgn46973;
    reg [31:0] z4697_assgn46974;
    reg [31:0] z4697_assgn46975;
    reg [31:0] z4697_assgn46976;
    reg [31:0] z1335_assgn1335;
    wire [31:0] b0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4701_assgn4701;
    reg [31:0] z4701_assgn47010;
    reg [31:0] z4701_assgn47011;
    reg [31:0] z4701_assgn47012;
    reg [31:0] z4701_assgn47013;
    reg [31:0] z4701_assgn47014;
    reg [31:0] z4701_assgn47015;
    reg [31:0] z4701_assgn47016;
    reg [31:0] z1337_assgn1337;
    wire [31:0] b1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4705_assgn4705;
    reg [31:0] z4705_assgn47050;
    reg [31:0] z4705_assgn47051;
    reg [31:0] z4705_assgn47052;
    reg [31:0] z4705_assgn47053;
    reg [31:0] z1339_assgn1339;
    reg [31:0] b0_G16_inv0_G256_inv0_reg;
    wire [31:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4709_assgn4709;
    reg [31:0] z4709_assgn47090;
    reg [31:0] z4709_assgn47091;
    reg [31:0] z4709_assgn47092;
    reg [31:0] z4709_assgn47093;
    reg [31:0] z1341_assgn1341;
    reg [31:0] b1_G16_inv0_G256_inv0_reg;
    wire [31:0] c1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4713_assgn4713;
    reg [31:0] z4713_assgn47130;
    reg [31:0] z4713_assgn47131;
    reg [31:0] z4713_assgn47132;
    reg [31:0] z4713_assgn47133;
    reg [31:0] z1343_assgn1343;
    wire [31:0] c0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4717_assgn4717;
    reg [31:0] z4717_assgn47170;
    reg [31:0] z4717_assgn47171;
    reg [31:0] z4717_assgn47172;
    reg [31:0] z4717_assgn47173;
    reg [31:0] z1345_assgn1345;
    wire [31:0] c1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4721_assgn4721;
    reg [31:0] z4721_assgn47210;
    reg [31:0] z4721_assgn47211;
    reg [31:0] z4721_assgn47212;
    reg [31:0] z4721_assgn47213;
    reg [31:0] z1347_assgn1347;
    wire [31:0] d0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4725_assgn4725;
    reg [31:0] z4725_assgn47250;
    reg [31:0] z4725_assgn47251;
    reg [31:0] z4725_assgn47252;
    reg [31:0] z4725_assgn47253;
    reg [31:0] z1349_assgn1349;
    wire [31:0] d1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] c0_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] d0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] axorb_1_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] c1_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] d1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4737_assgn4737;
    reg [31:0] z4737_assgn47370;
    reg [31:0] z4737_assgn47371;
    reg [31:0] z4737_assgn47372;
    reg [31:0] z4737_assgn47373;
    reg [31:0] z4737_assgn47374;
    reg [31:0] z1359_assgn1359;
    wire [31:0] r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4745_assgn4745;
    reg [31:0] z4745_assgn47450;
    reg [31:0] z1365_assgn1365;
    wire [31:0] u0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4749_assgn4749;
    reg [31:0] z4749_assgn47490;
    reg [31:0] z1367_assgn1367;
    wire [31:0] u1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] cxord_0_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] cxord_1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4757_assgn4757;
    reg [31:0] z4757_assgn47570;
    reg [31:0] z1373_assgn1373;
    wire [31:0] p0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] e0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4767_assgn4767;
    reg [31:0] z4767_assgn47670;
    reg [31:0] z1381_assgn1381;
    wire [31:0] p2_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] e1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4777_assgn4777;
    reg [31:0] z4777_assgn47770;
    reg [31:0] z4777_assgn47771;
    reg [31:0] z4777_assgn47772;
    reg [31:0] z4777_assgn47773;
    reg [31:0] z4777_assgn47774;
    reg [31:0] z1389_assgn1389;
    wire [31:0] r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4785_assgn4785;
    reg [31:0] z4785_assgn47850;
    reg [31:0] z1395_assgn1395;
    wire [31:0] u0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4789_assgn4789;
    reg [31:0] z4789_assgn47890;
    reg [31:0] z1397_assgn1397;
    wire [31:0] u1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4793_assgn4793;
    reg [31:0] z4793_assgn47930;
    reg [31:0] z1400_assgn1400;
    reg [31:0] r0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4797_assgn4797;
    reg [31:0] z4797_assgn47970;
    reg [31:0] z1402_assgn1402;
    wire [31:0] v1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4801_assgn4801;
    reg [31:0] z4801_assgn48010;
    reg [31:0] z4801_assgn48011;
    reg [31:0] z1403_assgn1403;
    wire [31:0] p0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4811_assgn4811;
    reg [31:0] z4811_assgn48110;
    reg [31:0] z4811_assgn48111;
    reg [31:0] z1411_assgn1411;
    wire [31:0] p2_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4825_assgn4825;
    reg [31:0] z4825_assgn48250;
    reg [31:0] z4825_assgn48251;
    reg [31:0] z4825_assgn48252;
    reg [31:0] z4825_assgn48253;
    reg [31:0] z4825_assgn48254;
    reg [31:0] z1423_assgn1423;
    wire [31:0] r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4833_assgn4833;
    reg [31:0] z4833_assgn48330;
    reg [31:0] z1429_assgn1429;
    wire [31:0] u0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4837_assgn4837;
    reg [31:0] z4837_assgn48370;
    reg [31:0] z1431_assgn1431;
    wire [31:0] u1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4841_assgn4841;
    reg [31:0] z4841_assgn48410;
    reg [31:0] z1434_assgn1434;
    reg [31:0] r0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4845_assgn4845;
    reg [31:0] z4845_assgn48450;
    reg [31:0] z1436_assgn1436;
    wire [31:0] v1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4849_assgn4849;
    reg [31:0] z4849_assgn48490;
    reg [31:0] z4849_assgn48491;
    reg [31:0] z1437_assgn1437;
    wire [31:0] p0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4859_assgn4859;
    reg [31:0] z4859_assgn48590;
    reg [31:0] z4859_assgn48591;
    reg [31:0] z1445_assgn1445;
    wire [31:0] p2_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4873_assgn4873;
    reg [31:0] z4873_assgn48730;
    reg [31:0] z4873_assgn48731;
    reg [31:0] z4873_assgn48732;
    reg [31:0] z4873_assgn48733;
    reg [31:0] z4873_assgn48734;
    reg [31:0] z4873_assgn48735;
    reg [31:0] z4873_assgn48736;
    reg [31:0] z4873_assgn48737;
    reg [31:0] z1457_assgn1457;
    wire [31:0] p1ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z4877_assgn4877;
    reg [31:0] z4877_assgn48770;
    reg [31:0] z4877_assgn48771;
    reg [31:0] z4877_assgn48772;
    reg [31:0] z4877_assgn48773;
    reg [31:0] z4877_assgn48774;
    reg [31:0] z4877_assgn48775;
    reg [31:0] z4877_assgn48776;
    reg [31:0] z4877_assgn48777;
    reg [31:0] z1459_assgn1459;
    wire [31:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p0_G16_inv0_G256_inv0;
    wire [31:0] p1_G16_inv0_G256_inv0;
    wire [31:0] z4885_assgn4885;
    reg [31:0] z4885_assgn48850;
    reg [31:0] z4885_assgn48851;
    reg [31:0] z4885_assgn48852;
    reg [31:0] z4885_assgn48853;
    reg [31:0] z1465_assgn1465;
    wire [31:0] r00_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4889_assgn4889;
    reg [31:0] z4889_assgn48890;
    reg [31:0] z4889_assgn48891;
    reg [31:0] z4889_assgn48892;
    reg [31:0] z4889_assgn48893;
    reg [31:0] z1467_assgn1467;
    wire [31:0] r10_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4893_assgn4893;
    reg [31:0] z4893_assgn48930;
    reg [31:0] z4893_assgn48931;
    reg [31:0] z4893_assgn48932;
    reg [31:0] z4893_assgn48933;
    reg [31:0] z1469_assgn1469;
    wire [31:0] r20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4897_assgn4897;
    reg [31:0] z4897_assgn48970;
    reg [31:0] z4897_assgn48971;
    reg [31:0] z4897_assgn48972;
    reg [31:0] z4897_assgn48973;
    reg [31:0] z4897_assgn48974;
    reg [31:0] z4897_assgn48975;
    reg [31:0] z4897_assgn48976;
    reg [31:0] z1471_assgn1471;
    wire [31:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4901_assgn4901;
    reg [31:0] z4901_assgn49010;
    reg [31:0] z4901_assgn49011;
    reg [31:0] z4901_assgn49012;
    reg [31:0] z4901_assgn49013;
    reg [31:0] z4901_assgn49014;
    reg [31:0] z4901_assgn49015;
    reg [31:0] z4901_assgn49016;
    reg [31:0] z1473_assgn1473;
    wire [31:0] a1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4905_assgn4905;
    reg [31:0] z4905_assgn49050;
    reg [31:0] z4905_assgn49051;
    reg [31:0] z4905_assgn49052;
    reg [31:0] z4905_assgn49053;
    reg [31:0] z4905_assgn49054;
    reg [31:0] z4905_assgn49055;
    reg [31:0] z4905_assgn49056;
    reg [31:0] z1475_assgn1475;
    wire [31:0] a0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4909_assgn4909;
    reg [31:0] z4909_assgn49090;
    reg [31:0] z4909_assgn49091;
    reg [31:0] z4909_assgn49092;
    reg [31:0] z4909_assgn49093;
    reg [31:0] z4909_assgn49094;
    reg [31:0] z4909_assgn49095;
    reg [31:0] z4909_assgn49096;
    reg [31:0] z1477_assgn1477;
    wire [31:0] a1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4913_assgn4913;
    reg [31:0] z4913_assgn49130;
    reg [31:0] z4913_assgn49131;
    reg [31:0] z4913_assgn49132;
    reg [31:0] z4913_assgn49133;
    reg [31:0] z4913_assgn49134;
    reg [31:0] z4913_assgn49135;
    reg [31:0] z4913_assgn49136;
    reg [31:0] z1479_assgn1479;
    wire [31:0] b0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4917_assgn4917;
    reg [31:0] z4917_assgn49170;
    reg [31:0] z4917_assgn49171;
    reg [31:0] z4917_assgn49172;
    reg [31:0] z4917_assgn49173;
    reg [31:0] z4917_assgn49174;
    reg [31:0] z4917_assgn49175;
    reg [31:0] z4917_assgn49176;
    reg [31:0] z1481_assgn1481;
    wire [31:0] b1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4921_assgn4921;
    reg [31:0] z4921_assgn49210;
    reg [31:0] z4921_assgn49211;
    reg [31:0] z4921_assgn49212;
    reg [31:0] z4921_assgn49213;
    reg [31:0] z1483_assgn1483;
    wire [31:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4925_assgn4925;
    reg [31:0] z4925_assgn49250;
    reg [31:0] z4925_assgn49251;
    reg [31:0] z4925_assgn49252;
    reg [31:0] z4925_assgn49253;
    reg [31:0] z1485_assgn1485;
    wire [31:0] c1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4929_assgn4929;
    reg [31:0] z4929_assgn49290;
    reg [31:0] z4929_assgn49291;
    reg [31:0] z4929_assgn49292;
    reg [31:0] z4929_assgn49293;
    reg [31:0] z1487_assgn1487;
    wire [31:0] c0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4933_assgn4933;
    reg [31:0] z4933_assgn49330;
    reg [31:0] z4933_assgn49331;
    reg [31:0] z4933_assgn49332;
    reg [31:0] z4933_assgn49333;
    reg [31:0] z1489_assgn1489;
    wire [31:0] c1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4937_assgn4937;
    reg [31:0] z4937_assgn49370;
    reg [31:0] z4937_assgn49371;
    reg [31:0] z4937_assgn49372;
    reg [31:0] z4937_assgn49373;
    reg [31:0] z1491_assgn1491;
    wire [31:0] d0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4941_assgn4941;
    reg [31:0] z4941_assgn49410;
    reg [31:0] z4941_assgn49411;
    reg [31:0] z4941_assgn49412;
    reg [31:0] z4941_assgn49413;
    reg [31:0] z1493_assgn1493;
    wire [31:0] d1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] c0_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] d0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] axorb_1_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] c1_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] d1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4953_assgn4953;
    reg [31:0] z4953_assgn49530;
    reg [31:0] z4953_assgn49531;
    reg [31:0] z4953_assgn49532;
    reg [31:0] z4953_assgn49533;
    reg [31:0] z4953_assgn49534;
    reg [31:0] z1503_assgn1503;
    wire [31:0] r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4961_assgn4961;
    reg [31:0] z4961_assgn49610;
    reg [31:0] z1509_assgn1509;
    wire [31:0] u0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4965_assgn4965;
    reg [31:0] z4965_assgn49650;
    reg [31:0] z1511_assgn1511;
    wire [31:0] u1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] cxord_0_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] cxord_1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4973_assgn4973;
    reg [31:0] z4973_assgn49730;
    reg [31:0] z1517_assgn1517;
    wire [31:0] p0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] e0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4983_assgn4983;
    reg [31:0] z4983_assgn49830;
    reg [31:0] z1525_assgn1525;
    wire [31:0] p2_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] e1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z4993_assgn4993;
    reg [31:0] z4993_assgn49930;
    reg [31:0] z4993_assgn49931;
    reg [31:0] z4993_assgn49932;
    reg [31:0] z4993_assgn49933;
    reg [31:0] z4993_assgn49934;
    reg [31:0] z1533_assgn1533;
    wire [31:0] r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5001_assgn5001;
    reg [31:0] z5001_assgn50010;
    reg [31:0] z1539_assgn1539;
    wire [31:0] u0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5005_assgn5005;
    reg [31:0] z5005_assgn50050;
    reg [31:0] z1541_assgn1541;
    wire [31:0] u1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5009_assgn5009;
    reg [31:0] z5009_assgn50090;
    reg [31:0] z1544_assgn1544;
    reg [31:0] r0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5013_assgn5013;
    reg [31:0] z5013_assgn50130;
    reg [31:0] z1546_assgn1546;
    wire [31:0] v1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5017_assgn5017;
    reg [31:0] z5017_assgn50170;
    reg [31:0] z5017_assgn50171;
    reg [31:0] z1547_assgn1547;
    wire [31:0] p0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5027_assgn5027;
    reg [31:0] z5027_assgn50270;
    reg [31:0] z5027_assgn50271;
    reg [31:0] z1555_assgn1555;
    wire [31:0] p2_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5041_assgn5041;
    reg [31:0] z5041_assgn50410;
    reg [31:0] z5041_assgn50411;
    reg [31:0] z5041_assgn50412;
    reg [31:0] z5041_assgn50413;
    reg [31:0] z5041_assgn50414;
    reg [31:0] z1567_assgn1567;
    wire [31:0] r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5049_assgn5049;
    reg [31:0] z5049_assgn50490;
    reg [31:0] z1573_assgn1573;
    wire [31:0] u0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5053_assgn5053;
    reg [31:0] z5053_assgn50530;
    reg [31:0] z1575_assgn1575;
    wire [31:0] u1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5057_assgn5057;
    reg [31:0] z5057_assgn50570;
    reg [31:0] z1578_assgn1578;
    reg [31:0] r0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5061_assgn5061;
    reg [31:0] z5061_assgn50610;
    reg [31:0] z1580_assgn1580;
    wire [31:0] v1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5065_assgn5065;
    reg [31:0] z5065_assgn50650;
    reg [31:0] z5065_assgn50651;
    reg [31:0] z1581_assgn1581;
    wire [31:0] p0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5075_assgn5075;
    reg [31:0] z5075_assgn50750;
    reg [31:0] z5075_assgn50751;
    reg [31:0] z1589_assgn1589;
    wire [31:0] p2_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5089_assgn5089;
    reg [31:0] z5089_assgn50890;
    reg [31:0] z5089_assgn50891;
    reg [31:0] z5089_assgn50892;
    reg [31:0] z5089_assgn50893;
    reg [31:0] z5089_assgn50894;
    reg [31:0] z5089_assgn50895;
    reg [31:0] z5089_assgn50896;
    reg [31:0] z5089_assgn50897;
    reg [31:0] z1601_assgn1601;
    wire [31:0] p1ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5093_assgn5093;
    reg [31:0] z5093_assgn50930;
    reg [31:0] z5093_assgn50931;
    reg [31:0] z5093_assgn50932;
    reg [31:0] z5093_assgn50933;
    reg [31:0] z5093_assgn50934;
    reg [31:0] z5093_assgn50935;
    reg [31:0] z5093_assgn50936;
    reg [31:0] z5093_assgn50937;
    reg [31:0] z1603_assgn1603;
    wire [31:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q0_G16_inv0_G256_inv0;
    wire [31:0] q1_G16_inv0_G256_inv0;
    wire [31:0] z5101_assgn5101;
    reg [31:0] z5101_assgn51010;
    reg [31:0] z5101_assgn51011;
    reg [31:0] z5101_assgn51012;
    reg [31:0] z5101_assgn51013;
    reg [31:0] z5101_assgn51014;
    reg [31:0] z5101_assgn51015;
    reg [31:0] z5101_assgn51016;
    reg [31:0] z5101_assgn51017;
    reg [31:0] z1609_assgn1609;
    wire [31:0] p0ls2_G16_inv0_G256_inv0;
    wire [31:0] z5105_assgn5105;
    reg [31:0] z5105_assgn51050;
    reg [31:0] z5105_assgn51051;
    reg [31:0] z5105_assgn51052;
    reg [31:0] z5105_assgn51053;
    reg [31:0] z5105_assgn51054;
    reg [31:0] z5105_assgn51055;
    reg [31:0] z5105_assgn51056;
    reg [31:0] z5105_assgn51057;
    reg [31:0] z1611_assgn1611;
    wire [31:0] p1ls2_G16_inv0_G256_inv0;
    wire [31:0] e0_G256_inv0;
    wire [31:0] e1_G256_inv0;
    wire [31:0] z5113_assgn5113;
    reg [31:0] z5113_assgn51130;
    reg [31:0] z5113_assgn51131;
    reg [31:0] z5113_assgn51132;
    reg [31:0] z5113_assgn51133;
    reg [31:0] z5113_assgn51134;
    reg [31:0] z1617_assgn1617;
    wire [31:0] r00_G16_mul1_G256_inv0;
    wire [31:0] z5117_assgn5117;
    reg [31:0] z5117_assgn51170;
    reg [31:0] z5117_assgn51171;
    reg [31:0] z5117_assgn51172;
    reg [31:0] z5117_assgn51173;
    reg [31:0] z5117_assgn51174;
    reg [31:0] z1619_assgn1619;
    wire [31:0] r10_G16_mul1_G256_inv0;
    wire [31:0] z5121_assgn5121;
    reg [31:0] z5121_assgn51210;
    reg [31:0] z5121_assgn51211;
    reg [31:0] z5121_assgn51212;
    reg [31:0] z5121_assgn51213;
    reg [31:0] z5121_assgn51214;
    reg [31:0] z1621_assgn1621;
    wire [31:0] r20_G16_mul1_G256_inv0;
    wire [31:0] z5125_assgn5125;
    reg [31:0] z5125_assgn51250;
    reg [31:0] z5125_assgn51251;
    reg [31:0] z5125_assgn51252;
    reg [31:0] z5125_assgn51253;
    reg [31:0] z5125_assgn51254;
    reg [31:0] z1623_assgn1623;
    wire [31:0] r30_G16_mul1_G256_inv0;
    wire [31:0] z5129_assgn5129;
    reg [31:0] z5129_assgn51290;
    reg [31:0] z5129_assgn51291;
    reg [31:0] z5129_assgn51292;
    reg [31:0] z5129_assgn51293;
    reg [31:0] z5129_assgn51294;
    reg [31:0] z1625_assgn1625;
    wire [31:0] r40_G16_mul1_G256_inv0;
    wire [31:0] z5133_assgn5133;
    reg [31:0] z5133_assgn51330;
    reg [31:0] z5133_assgn51331;
    reg [31:0] z5133_assgn51332;
    reg [31:0] z5133_assgn51333;
    reg [31:0] z5133_assgn51334;
    reg [31:0] z1627_assgn1627;
    wire [31:0] r50_G16_mul1_G256_inv0;
    wire [31:0] z5137_assgn5137;
    reg [31:0] z5137_assgn51370;
    reg [31:0] z5137_assgn51371;
    reg [31:0] z5137_assgn51372;
    reg [31:0] z5137_assgn51373;
    reg [31:0] z5137_assgn51374;
    reg [31:0] z1629_assgn1629;
    wire [31:0] r60_G16_mul1_G256_inv0;
    wire [31:0] z5141_assgn5141;
    reg [31:0] z5141_assgn51410;
    reg [31:0] z5141_assgn51411;
    reg [31:0] z5141_assgn51412;
    reg [31:0] z5141_assgn51413;
    reg [31:0] z5141_assgn51414;
    reg [31:0] z1631_assgn1631;
    wire [31:0] r70_G16_mul1_G256_inv0;
    wire [31:0] z5145_assgn5145;
    reg [31:0] z5145_assgn51450;
    reg [31:0] z5145_assgn51451;
    reg [31:0] z5145_assgn51452;
    reg [31:0] z5145_assgn51453;
    reg [31:0] z5145_assgn51454;
    reg [31:0] z1633_assgn1633;
    wire [31:0] r80_G16_mul1_G256_inv0;
    wire [31:0] z5149_assgn5149;
    reg [31:0] z5149_assgn51490;
    reg [31:0] z5149_assgn51491;
    reg [31:0] z5149_assgn51492;
    reg [31:0] z5149_assgn51493;
    reg [31:0] z5149_assgn51494;
    reg [31:0] z5149_assgn51495;
    reg [31:0] z5149_assgn51496;
    reg [31:0] z5149_assgn51497;
    reg [31:0] z1635_assgn1635;
    wire [31:0] a0_0_G16_mul1_G256_inv0;
    wire [31:0] z5153_assgn5153;
    reg [31:0] z5153_assgn51530;
    reg [31:0] z5153_assgn51531;
    reg [31:0] z5153_assgn51532;
    reg [31:0] z5153_assgn51533;
    reg [31:0] z5153_assgn51534;
    reg [31:0] z5153_assgn51535;
    reg [31:0] z5153_assgn51536;
    reg [31:0] z5153_assgn51537;
    reg [31:0] z1637_assgn1637;
    wire [31:0] a1_0_G16_mul1_G256_inv0;
    wire [31:0] z5157_assgn5157;
    reg [31:0] z5157_assgn51570;
    reg [31:0] z5157_assgn51571;
    reg [31:0] z5157_assgn51572;
    reg [31:0] z5157_assgn51573;
    reg [31:0] z5157_assgn51574;
    reg [31:0] z5157_assgn51575;
    reg [31:0] z5157_assgn51576;
    reg [31:0] z5157_assgn51577;
    reg [31:0] z1639_assgn1639;
    wire [31:0] a0_G16_mul1_G256_inv0;
    wire [31:0] z5161_assgn5161;
    reg [31:0] z5161_assgn51610;
    reg [31:0] z5161_assgn51611;
    reg [31:0] z5161_assgn51612;
    reg [31:0] z5161_assgn51613;
    reg [31:0] z5161_assgn51614;
    reg [31:0] z5161_assgn51615;
    reg [31:0] z5161_assgn51616;
    reg [31:0] z5161_assgn51617;
    reg [31:0] z1641_assgn1641;
    wire [31:0] a1_G16_mul1_G256_inv0;
    wire [31:0] z5165_assgn5165;
    reg [31:0] z5165_assgn51650;
    reg [31:0] z5165_assgn51651;
    reg [31:0] z5165_assgn51652;
    reg [31:0] z5165_assgn51653;
    reg [31:0] z5165_assgn51654;
    reg [31:0] z5165_assgn51655;
    reg [31:0] z5165_assgn51656;
    reg [31:0] z5165_assgn51657;
    reg [31:0] z1643_assgn1643;
    wire [31:0] b0_G16_mul1_G256_inv0;
    wire [31:0] z5169_assgn5169;
    reg [31:0] z5169_assgn51690;
    reg [31:0] z5169_assgn51691;
    reg [31:0] z5169_assgn51692;
    reg [31:0] z5169_assgn51693;
    reg [31:0] z5169_assgn51694;
    reg [31:0] z5169_assgn51695;
    reg [31:0] z5169_assgn51696;
    reg [31:0] z5169_assgn51697;
    reg [31:0] z1645_assgn1645;
    wire [31:0] b1_G16_mul1_G256_inv0;
    wire [31:0] z5173_assgn5173;
    reg [31:0] z5173_assgn51730;
    reg [31:0] z5173_assgn51731;
    reg [31:0] z5173_assgn51732;
    reg [31:0] z5173_assgn51733;
    reg [31:0] z5173_assgn51734;
    reg [31:0] z1647_assgn1647;
    wire [31:0] z5175_assgn5175;
    reg [31:0] z5175_assgn51750;
    reg [31:0] z5175_assgn51751;
    reg [31:0] z5175_assgn51752;
    reg [31:0] z5175_assgn51753;
    reg [31:0] z5175_assgn51754;
    reg [31:0] z1648_assgn1648;
    wire [31:0] c0_0_G16_mul1_G256_inv0;
    wire [31:0] z5179_assgn5179;
    reg [31:0] z5179_assgn51790;
    reg [31:0] z5179_assgn51791;
    reg [31:0] z5179_assgn51792;
    reg [31:0] z5179_assgn51793;
    reg [31:0] z5179_assgn51794;
    reg [31:0] z1649_assgn1649;
    wire [31:0] z5181_assgn5181;
    reg [31:0] z5181_assgn51810;
    reg [31:0] z5181_assgn51811;
    reg [31:0] z5181_assgn51812;
    reg [31:0] z5181_assgn51813;
    reg [31:0] z5181_assgn51814;
    reg [31:0] z1650_assgn1650;
    wire [31:0] c1_0_G16_mul1_G256_inv0;
    wire [31:0] z5185_assgn5185;
    reg [31:0] z5185_assgn51850;
    reg [31:0] z5185_assgn51851;
    reg [31:0] z5185_assgn51852;
    reg [31:0] z5185_assgn51853;
    reg [31:0] z5185_assgn51854;
    reg [31:0] z1651_assgn1651;
    wire [31:0] c0_G16_mul1_G256_inv0;
    wire [31:0] z5189_assgn5189;
    reg [31:0] z5189_assgn51890;
    reg [31:0] z5189_assgn51891;
    reg [31:0] z5189_assgn51892;
    reg [31:0] z5189_assgn51893;
    reg [31:0] z5189_assgn51894;
    reg [31:0] z1653_assgn1653;
    wire [31:0] c1_G16_mul1_G256_inv0;
    wire [31:0] z5193_assgn5193;
    reg [31:0] z5193_assgn51930;
    reg [31:0] z5193_assgn51931;
    reg [31:0] z5193_assgn51932;
    reg [31:0] z5193_assgn51933;
    reg [31:0] z5193_assgn51934;
    reg [31:0] z1655_assgn1655;
    wire [31:0] z5195_assgn5195;
    reg [31:0] z5195_assgn51950;
    reg [31:0] z5195_assgn51951;
    reg [31:0] z5195_assgn51952;
    reg [31:0] z5195_assgn51953;
    reg [31:0] z5195_assgn51954;
    reg [31:0] z1656_assgn1656;
    wire [31:0] d0_G16_mul1_G256_inv0;
    wire [31:0] z5199_assgn5199;
    reg [31:0] z5199_assgn51990;
    reg [31:0] z5199_assgn51991;
    reg [31:0] z5199_assgn51992;
    reg [31:0] z5199_assgn51993;
    reg [31:0] z5199_assgn51994;
    reg [31:0] z1657_assgn1657;
    wire [31:0] z5201_assgn5201;
    reg [31:0] z5201_assgn52010;
    reg [31:0] z5201_assgn52011;
    reg [31:0] z5201_assgn52012;
    reg [31:0] z5201_assgn52013;
    reg [31:0] z5201_assgn52014;
    reg [31:0] z1658_assgn1658;
    wire [31:0] d1_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G16_mul1_G256_inv0;
    wire [31:0] cxord_0_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G16_mul1_G256_inv0;
    wire [31:0] cxord_1_G16_mul1_G256_inv0;
    wire [31:0] z5213_assgn5213;
    reg [31:0] z5213_assgn52130;
    reg [31:0] z5213_assgn52131;
    reg [31:0] z5213_assgn52132;
    reg [31:0] z5213_assgn52133;
    reg [31:0] z5213_assgn52134;
    reg [31:0] z1667_assgn1667;
    wire [31:0] r00_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5217_assgn5217;
    reg [31:0] z5217_assgn52170;
    reg [31:0] z5217_assgn52171;
    reg [31:0] z5217_assgn52172;
    reg [31:0] z5217_assgn52173;
    reg [31:0] z5217_assgn52174;
    reg [31:0] z1669_assgn1669;
    wire [31:0] r10_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5221_assgn5221;
    reg [31:0] z5221_assgn52210;
    reg [31:0] z5221_assgn52211;
    reg [31:0] z5221_assgn52212;
    reg [31:0] z5221_assgn52213;
    reg [31:0] z5221_assgn52214;
    reg [31:0] z1671_assgn1671;
    wire [31:0] r20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5225_assgn5225;
    reg [31:0] z5225_assgn52250;
    reg [31:0] z5225_assgn52251;
    reg [31:0] z5225_assgn52252;
    reg [31:0] z5225_assgn52253;
    reg [31:0] z5225_assgn52254;
    reg [31:0] z5225_assgn52255;
    reg [31:0] z5225_assgn52256;
    reg [31:0] z5225_assgn52257;
    reg [31:0] z1673_assgn1673;
    wire [31:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5229_assgn5229;
    reg [31:0] z5229_assgn52290;
    reg [31:0] z5229_assgn52291;
    reg [31:0] z5229_assgn52292;
    reg [31:0] z5229_assgn52293;
    reg [31:0] z5229_assgn52294;
    reg [31:0] z5229_assgn52295;
    reg [31:0] z5229_assgn52296;
    reg [31:0] z5229_assgn52297;
    reg [31:0] z1675_assgn1675;
    wire [31:0] a1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5233_assgn5233;
    reg [31:0] z5233_assgn52330;
    reg [31:0] z5233_assgn52331;
    reg [31:0] z5233_assgn52332;
    reg [31:0] z5233_assgn52333;
    reg [31:0] z5233_assgn52334;
    reg [31:0] z5233_assgn52335;
    reg [31:0] z5233_assgn52336;
    reg [31:0] z5233_assgn52337;
    reg [31:0] z1677_assgn1677;
    wire [31:0] a0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5237_assgn5237;
    reg [31:0] z5237_assgn52370;
    reg [31:0] z5237_assgn52371;
    reg [31:0] z5237_assgn52372;
    reg [31:0] z5237_assgn52373;
    reg [31:0] z5237_assgn52374;
    reg [31:0] z5237_assgn52375;
    reg [31:0] z5237_assgn52376;
    reg [31:0] z5237_assgn52377;
    reg [31:0] z1679_assgn1679;
    wire [31:0] a1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5241_assgn5241;
    reg [31:0] z5241_assgn52410;
    reg [31:0] z5241_assgn52411;
    reg [31:0] z5241_assgn52412;
    reg [31:0] z5241_assgn52413;
    reg [31:0] z5241_assgn52414;
    reg [31:0] z5241_assgn52415;
    reg [31:0] z5241_assgn52416;
    reg [31:0] z5241_assgn52417;
    reg [31:0] z1681_assgn1681;
    wire [31:0] b0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5245_assgn5245;
    reg [31:0] z5245_assgn52450;
    reg [31:0] z5245_assgn52451;
    reg [31:0] z5245_assgn52452;
    reg [31:0] z5245_assgn52453;
    reg [31:0] z5245_assgn52454;
    reg [31:0] z5245_assgn52455;
    reg [31:0] z5245_assgn52456;
    reg [31:0] z5245_assgn52457;
    reg [31:0] z1683_assgn1683;
    wire [31:0] b1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5249_assgn5249;
    reg [31:0] z5249_assgn52490;
    reg [31:0] z5249_assgn52491;
    reg [31:0] z5249_assgn52492;
    reg [31:0] z5249_assgn52493;
    reg [31:0] z5249_assgn52494;
    reg [31:0] z1685_assgn1685;
    wire [31:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5253_assgn5253;
    reg [31:0] z5253_assgn52530;
    reg [31:0] z5253_assgn52531;
    reg [31:0] z5253_assgn52532;
    reg [31:0] z5253_assgn52533;
    reg [31:0] z5253_assgn52534;
    reg [31:0] z1687_assgn1687;
    wire [31:0] c1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5257_assgn5257;
    reg [31:0] z5257_assgn52570;
    reg [31:0] z5257_assgn52571;
    reg [31:0] z5257_assgn52572;
    reg [31:0] z5257_assgn52573;
    reg [31:0] z5257_assgn52574;
    reg [31:0] z1689_assgn1689;
    wire [31:0] c0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5261_assgn5261;
    reg [31:0] z5261_assgn52610;
    reg [31:0] z5261_assgn52611;
    reg [31:0] z5261_assgn52612;
    reg [31:0] z5261_assgn52613;
    reg [31:0] z5261_assgn52614;
    reg [31:0] z1691_assgn1691;
    wire [31:0] c1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5265_assgn5265;
    reg [31:0] z5265_assgn52650;
    reg [31:0] z5265_assgn52651;
    reg [31:0] z5265_assgn52652;
    reg [31:0] z5265_assgn52653;
    reg [31:0] z5265_assgn52654;
    reg [31:0] z1693_assgn1693;
    wire [31:0] d0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5269_assgn5269;
    reg [31:0] z5269_assgn52690;
    reg [31:0] z5269_assgn52691;
    reg [31:0] z5269_assgn52692;
    reg [31:0] z5269_assgn52693;
    reg [31:0] z5269_assgn52694;
    reg [31:0] z1695_assgn1695;
    wire [31:0] d1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] c0_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] d0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] c1_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] d1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5281_assgn5281;
    reg [31:0] z5281_assgn52810;
    reg [31:0] z5281_assgn52811;
    reg [31:0] z5281_assgn52812;
    reg [31:0] z5281_assgn52813;
    reg [31:0] z5281_assgn52814;
    reg [31:0] z5281_assgn52815;
    reg [31:0] z1705_assgn1705;
    wire [31:0] r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5289_assgn5289;
    reg [31:0] z5289_assgn52890;
    reg [31:0] z1711_assgn1711;
    wire [31:0] u0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5293_assgn5293;
    reg [31:0] z5293_assgn52930;
    reg [31:0] z1713_assgn1713;
    wire [31:0] u1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] cxord_0_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] cxord_1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5301_assgn5301;
    reg [31:0] z5301_assgn53010;
    reg [31:0] z1719_assgn1719;
    wire [31:0] p0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] e0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5311_assgn5311;
    reg [31:0] z5311_assgn53110;
    reg [31:0] z1727_assgn1727;
    wire [31:0] p2_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] e1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5321_assgn5321;
    reg [31:0] z5321_assgn53210;
    reg [31:0] z5321_assgn53211;
    reg [31:0] z5321_assgn53212;
    reg [31:0] z5321_assgn53213;
    reg [31:0] z5321_assgn53214;
    reg [31:0] z5321_assgn53215;
    reg [31:0] z1735_assgn1735;
    wire [31:0] r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5329_assgn5329;
    reg [31:0] z5329_assgn53290;
    reg [31:0] z1741_assgn1741;
    wire [31:0] u0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5333_assgn5333;
    reg [31:0] z5333_assgn53330;
    reg [31:0] z1743_assgn1743;
    wire [31:0] u1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5337_assgn5337;
    reg [31:0] z5337_assgn53370;
    reg [31:0] z1746_assgn1746;
    reg [31:0] r0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5341_assgn5341;
    reg [31:0] z5341_assgn53410;
    reg [31:0] z1748_assgn1748;
    wire [31:0] v1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5345_assgn5345;
    reg [31:0] z5345_assgn53450;
    reg [31:0] z5345_assgn53451;
    reg [31:0] z1749_assgn1749;
    wire [31:0] p0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5355_assgn5355;
    reg [31:0] z5355_assgn53550;
    reg [31:0] z5355_assgn53551;
    reg [31:0] z1757_assgn1757;
    wire [31:0] p2_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5369_assgn5369;
    reg [31:0] z5369_assgn53690;
    reg [31:0] z5369_assgn53691;
    reg [31:0] z5369_assgn53692;
    reg [31:0] z5369_assgn53693;
    reg [31:0] z5369_assgn53694;
    reg [31:0] z5369_assgn53695;
    reg [31:0] z1769_assgn1769;
    wire [31:0] r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5377_assgn5377;
    reg [31:0] z5377_assgn53770;
    reg [31:0] z1775_assgn1775;
    wire [31:0] u0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5381_assgn5381;
    reg [31:0] z5381_assgn53810;
    reg [31:0] z1777_assgn1777;
    wire [31:0] u1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5385_assgn5385;
    reg [31:0] z5385_assgn53850;
    reg [31:0] z1780_assgn1780;
    reg [31:0] r0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5389_assgn5389;
    reg [31:0] z5389_assgn53890;
    reg [31:0] z1782_assgn1782;
    wire [31:0] v1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5393_assgn5393;
    reg [31:0] z5393_assgn53930;
    reg [31:0] z5393_assgn53931;
    reg [31:0] z1783_assgn1783;
    wire [31:0] p0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5403_assgn5403;
    reg [31:0] z5403_assgn54030;
    reg [31:0] z5403_assgn54031;
    reg [31:0] z1791_assgn1791;
    wire [31:0] p2_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5417_assgn5417;
    reg [31:0] z5417_assgn54170;
    reg [31:0] z5417_assgn54171;
    reg [31:0] z5417_assgn54172;
    reg [31:0] z5417_assgn54173;
    reg [31:0] z5417_assgn54174;
    reg [31:0] z5417_assgn54175;
    reg [31:0] z5417_assgn54176;
    reg [31:0] z5417_assgn54177;
    reg [31:0] z5417_assgn54178;
    reg [31:0] z1803_assgn1803;
    wire [31:0] p1ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5421_assgn5421;
    reg [31:0] z5421_assgn54210;
    reg [31:0] z5421_assgn54211;
    reg [31:0] z5421_assgn54212;
    reg [31:0] z5421_assgn54213;
    reg [31:0] z5421_assgn54214;
    reg [31:0] z5421_assgn54215;
    reg [31:0] z5421_assgn54216;
    reg [31:0] z5421_assgn54217;
    reg [31:0] z5421_assgn54218;
    reg [31:0] z1805_assgn1805;
    wire [31:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] e0_G16_mul1_G256_inv0;
    wire [31:0] e1_G16_mul1_G256_inv0;
    wire [31:0] z5429_assgn5429;
    reg [31:0] z5429_assgn54290;
    reg [31:0] z5429_assgn54291;
    reg [31:0] z5429_assgn54292;
    reg [31:0] z5429_assgn54293;
    reg [31:0] z5429_assgn54294;
    reg [31:0] z5429_assgn54295;
    reg [31:0] z5429_assgn54296;
    reg [31:0] z5429_assgn54297;
    reg [31:0] z5429_assgn54298;
    reg [31:0] z1811_assgn1811;
    wire [31:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5433_assgn5433;
    reg [31:0] z5433_assgn54330;
    reg [31:0] z5433_assgn54331;
    reg [31:0] z5433_assgn54332;
    reg [31:0] z5433_assgn54333;
    reg [31:0] z5433_assgn54334;
    reg [31:0] z5433_assgn54335;
    reg [31:0] z5433_assgn54336;
    reg [31:0] z5433_assgn54337;
    reg [31:0] z5433_assgn54338;
    reg [31:0] z1813_assgn1813;
    wire [31:0] a1_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5437_assgn5437;
    reg [31:0] z5437_assgn54370;
    reg [31:0] z5437_assgn54371;
    reg [31:0] z5437_assgn54372;
    reg [31:0] z5437_assgn54373;
    reg [31:0] z5437_assgn54374;
    reg [31:0] z5437_assgn54375;
    reg [31:0] z5437_assgn54376;
    reg [31:0] z5437_assgn54377;
    reg [31:0] z5437_assgn54378;
    reg [31:0] z1815_assgn1815;
    wire [31:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5441_assgn5441;
    reg [31:0] z5441_assgn54410;
    reg [31:0] z5441_assgn54411;
    reg [31:0] z5441_assgn54412;
    reg [31:0] z5441_assgn54413;
    reg [31:0] z5441_assgn54414;
    reg [31:0] z5441_assgn54415;
    reg [31:0] z5441_assgn54416;
    reg [31:0] z5441_assgn54417;
    reg [31:0] z5441_assgn54418;
    reg [31:0] z1817_assgn1817;
    wire [31:0] a1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5445_assgn5445;
    reg [31:0] z5445_assgn54450;
    reg [31:0] z5445_assgn54451;
    reg [31:0] z5445_assgn54452;
    reg [31:0] z5445_assgn54453;
    reg [31:0] z5445_assgn54454;
    reg [31:0] z5445_assgn54455;
    reg [31:0] z5445_assgn54456;
    reg [31:0] z5445_assgn54457;
    reg [31:0] z5445_assgn54458;
    reg [31:0] z1819_assgn1819;
    wire [31:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5449_assgn5449;
    reg [31:0] z5449_assgn54490;
    reg [31:0] z5449_assgn54491;
    reg [31:0] z5449_assgn54492;
    reg [31:0] z5449_assgn54493;
    reg [31:0] z5449_assgn54494;
    reg [31:0] z5449_assgn54495;
    reg [31:0] z5449_assgn54496;
    reg [31:0] z5449_assgn54497;
    reg [31:0] z5449_assgn54498;
    reg [31:0] z1821_assgn1821;
    wire [31:0] b1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5461_assgn5461;
    reg [31:0] z5461_assgn54610;
    reg [31:0] z5461_assgn54611;
    reg [31:0] z5461_assgn54612;
    reg [31:0] z5461_assgn54613;
    reg [31:0] z5461_assgn54614;
    reg [31:0] z5461_assgn54615;
    reg [31:0] z5461_assgn54616;
    reg [31:0] z5461_assgn54617;
    reg [31:0] z5461_assgn54618;
    reg [31:0] z1831_assgn1831;
    wire [31:0] p1ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z5465_assgn5465;
    reg [31:0] z5465_assgn54650;
    reg [31:0] z5465_assgn54651;
    reg [31:0] z5465_assgn54652;
    reg [31:0] z5465_assgn54653;
    reg [31:0] z5465_assgn54654;
    reg [31:0] z5465_assgn54655;
    reg [31:0] z5465_assgn54656;
    reg [31:0] z5465_assgn54657;
    reg [31:0] z5465_assgn54658;
    reg [31:0] z1833_assgn1833;
    wire [31:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] e01_G16_mul1_G256_inv0;
    wire [31:0] e11_G16_mul1_G256_inv0;
    wire [31:0] z5473_assgn5473;
    reg [31:0] z5473_assgn54730;
    reg [31:0] z5473_assgn54731;
    reg [31:0] z5473_assgn54732;
    reg [31:0] z5473_assgn54733;
    reg [31:0] z5473_assgn54734;
    reg [31:0] z1839_assgn1839;
    wire [31:0] r00_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5477_assgn5477;
    reg [31:0] z5477_assgn54770;
    reg [31:0] z5477_assgn54771;
    reg [31:0] z5477_assgn54772;
    reg [31:0] z5477_assgn54773;
    reg [31:0] z5477_assgn54774;
    reg [31:0] z1841_assgn1841;
    wire [31:0] r10_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5481_assgn5481;
    reg [31:0] z5481_assgn54810;
    reg [31:0] z5481_assgn54811;
    reg [31:0] z5481_assgn54812;
    reg [31:0] z5481_assgn54813;
    reg [31:0] z5481_assgn54814;
    reg [31:0] z1843_assgn1843;
    wire [31:0] r20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5485_assgn5485;
    reg [31:0] z5485_assgn54850;
    reg [31:0] z5485_assgn54851;
    reg [31:0] z5485_assgn54852;
    reg [31:0] z5485_assgn54853;
    reg [31:0] z5485_assgn54854;
    reg [31:0] z5485_assgn54855;
    reg [31:0] z5485_assgn54856;
    reg [31:0] z5485_assgn54857;
    reg [31:0] z1845_assgn1845;
    wire [31:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5489_assgn5489;
    reg [31:0] z5489_assgn54890;
    reg [31:0] z5489_assgn54891;
    reg [31:0] z5489_assgn54892;
    reg [31:0] z5489_assgn54893;
    reg [31:0] z5489_assgn54894;
    reg [31:0] z5489_assgn54895;
    reg [31:0] z5489_assgn54896;
    reg [31:0] z5489_assgn54897;
    reg [31:0] z1847_assgn1847;
    wire [31:0] a1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5493_assgn5493;
    reg [31:0] z5493_assgn54930;
    reg [31:0] z5493_assgn54931;
    reg [31:0] z5493_assgn54932;
    reg [31:0] z5493_assgn54933;
    reg [31:0] z5493_assgn54934;
    reg [31:0] z5493_assgn54935;
    reg [31:0] z5493_assgn54936;
    reg [31:0] z5493_assgn54937;
    reg [31:0] z1849_assgn1849;
    wire [31:0] a0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5497_assgn5497;
    reg [31:0] z5497_assgn54970;
    reg [31:0] z5497_assgn54971;
    reg [31:0] z5497_assgn54972;
    reg [31:0] z5497_assgn54973;
    reg [31:0] z5497_assgn54974;
    reg [31:0] z5497_assgn54975;
    reg [31:0] z5497_assgn54976;
    reg [31:0] z5497_assgn54977;
    reg [31:0] z1851_assgn1851;
    wire [31:0] a1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5501_assgn5501;
    reg [31:0] z5501_assgn55010;
    reg [31:0] z5501_assgn55011;
    reg [31:0] z5501_assgn55012;
    reg [31:0] z5501_assgn55013;
    reg [31:0] z5501_assgn55014;
    reg [31:0] z5501_assgn55015;
    reg [31:0] z5501_assgn55016;
    reg [31:0] z5501_assgn55017;
    reg [31:0] z1853_assgn1853;
    wire [31:0] b0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5505_assgn5505;
    reg [31:0] z5505_assgn55050;
    reg [31:0] z5505_assgn55051;
    reg [31:0] z5505_assgn55052;
    reg [31:0] z5505_assgn55053;
    reg [31:0] z5505_assgn55054;
    reg [31:0] z5505_assgn55055;
    reg [31:0] z5505_assgn55056;
    reg [31:0] z5505_assgn55057;
    reg [31:0] z1855_assgn1855;
    wire [31:0] b1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5509_assgn5509;
    reg [31:0] z5509_assgn55090;
    reg [31:0] z5509_assgn55091;
    reg [31:0] z5509_assgn55092;
    reg [31:0] z5509_assgn55093;
    reg [31:0] z5509_assgn55094;
    reg [31:0] z1857_assgn1857;
    wire [31:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5513_assgn5513;
    reg [31:0] z5513_assgn55130;
    reg [31:0] z5513_assgn55131;
    reg [31:0] z5513_assgn55132;
    reg [31:0] z5513_assgn55133;
    reg [31:0] z5513_assgn55134;
    reg [31:0] z1859_assgn1859;
    wire [31:0] c1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5517_assgn5517;
    reg [31:0] z5517_assgn55170;
    reg [31:0] z5517_assgn55171;
    reg [31:0] z5517_assgn55172;
    reg [31:0] z5517_assgn55173;
    reg [31:0] z5517_assgn55174;
    reg [31:0] z1861_assgn1861;
    wire [31:0] c0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5521_assgn5521;
    reg [31:0] z5521_assgn55210;
    reg [31:0] z5521_assgn55211;
    reg [31:0] z5521_assgn55212;
    reg [31:0] z5521_assgn55213;
    reg [31:0] z5521_assgn55214;
    reg [31:0] z1863_assgn1863;
    wire [31:0] c1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5525_assgn5525;
    reg [31:0] z5525_assgn55250;
    reg [31:0] z5525_assgn55251;
    reg [31:0] z5525_assgn55252;
    reg [31:0] z5525_assgn55253;
    reg [31:0] z5525_assgn55254;
    reg [31:0] z1865_assgn1865;
    wire [31:0] d0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5529_assgn5529;
    reg [31:0] z5529_assgn55290;
    reg [31:0] z5529_assgn55291;
    reg [31:0] z5529_assgn55292;
    reg [31:0] z5529_assgn55293;
    reg [31:0] z5529_assgn55294;
    reg [31:0] z1867_assgn1867;
    wire [31:0] d1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] c0_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] d0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] c1_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] d1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5541_assgn5541;
    reg [31:0] z5541_assgn55410;
    reg [31:0] z5541_assgn55411;
    reg [31:0] z5541_assgn55412;
    reg [31:0] z5541_assgn55413;
    reg [31:0] z5541_assgn55414;
    reg [31:0] z5541_assgn55415;
    reg [31:0] z1877_assgn1877;
    wire [31:0] r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5549_assgn5549;
    reg [31:0] z5549_assgn55490;
    reg [31:0] z1883_assgn1883;
    wire [31:0] u0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5553_assgn5553;
    reg [31:0] z5553_assgn55530;
    reg [31:0] z1885_assgn1885;
    wire [31:0] u1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] cxord_0_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] cxord_1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5561_assgn5561;
    reg [31:0] z5561_assgn55610;
    reg [31:0] z1891_assgn1891;
    wire [31:0] p0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] e0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5571_assgn5571;
    reg [31:0] z5571_assgn55710;
    reg [31:0] z1899_assgn1899;
    wire [31:0] p2_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] e1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5581_assgn5581;
    reg [31:0] z5581_assgn55810;
    reg [31:0] z5581_assgn55811;
    reg [31:0] z5581_assgn55812;
    reg [31:0] z5581_assgn55813;
    reg [31:0] z5581_assgn55814;
    reg [31:0] z5581_assgn55815;
    reg [31:0] z1907_assgn1907;
    wire [31:0] r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5589_assgn5589;
    reg [31:0] z5589_assgn55890;
    reg [31:0] z1913_assgn1913;
    wire [31:0] u0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5593_assgn5593;
    reg [31:0] z5593_assgn55930;
    reg [31:0] z1915_assgn1915;
    wire [31:0] u1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5597_assgn5597;
    reg [31:0] z5597_assgn55970;
    reg [31:0] z1918_assgn1918;
    reg [31:0] r0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5601_assgn5601;
    reg [31:0] z5601_assgn56010;
    reg [31:0] z1920_assgn1920;
    wire [31:0] v1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5605_assgn5605;
    reg [31:0] z5605_assgn56050;
    reg [31:0] z5605_assgn56051;
    reg [31:0] z1921_assgn1921;
    wire [31:0] p0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5615_assgn5615;
    reg [31:0] z5615_assgn56150;
    reg [31:0] z5615_assgn56151;
    reg [31:0] z1929_assgn1929;
    wire [31:0] p2_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5629_assgn5629;
    reg [31:0] z5629_assgn56290;
    reg [31:0] z5629_assgn56291;
    reg [31:0] z5629_assgn56292;
    reg [31:0] z5629_assgn56293;
    reg [31:0] z5629_assgn56294;
    reg [31:0] z5629_assgn56295;
    reg [31:0] z1941_assgn1941;
    wire [31:0] r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5637_assgn5637;
    reg [31:0] z5637_assgn56370;
    reg [31:0] z1947_assgn1947;
    wire [31:0] u0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5641_assgn5641;
    reg [31:0] z5641_assgn56410;
    reg [31:0] z1949_assgn1949;
    wire [31:0] u1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5645_assgn5645;
    reg [31:0] z5645_assgn56450;
    reg [31:0] z1952_assgn1952;
    reg [31:0] r0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5649_assgn5649;
    reg [31:0] z5649_assgn56490;
    reg [31:0] z1954_assgn1954;
    wire [31:0] v1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5653_assgn5653;
    reg [31:0] z5653_assgn56530;
    reg [31:0] z5653_assgn56531;
    reg [31:0] z1955_assgn1955;
    wire [31:0] p0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5663_assgn5663;
    reg [31:0] z5663_assgn56630;
    reg [31:0] z5663_assgn56631;
    reg [31:0] z1963_assgn1963;
    wire [31:0] p2_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5677_assgn5677;
    reg [31:0] z5677_assgn56770;
    reg [31:0] z5677_assgn56771;
    reg [31:0] z5677_assgn56772;
    reg [31:0] z5677_assgn56773;
    reg [31:0] z5677_assgn56774;
    reg [31:0] z5677_assgn56775;
    reg [31:0] z5677_assgn56776;
    reg [31:0] z5677_assgn56777;
    reg [31:0] z5677_assgn56778;
    reg [31:0] z1975_assgn1975;
    wire [31:0] p1ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z5681_assgn5681;
    reg [31:0] z5681_assgn56810;
    reg [31:0] z5681_assgn56811;
    reg [31:0] z5681_assgn56812;
    reg [31:0] z5681_assgn56813;
    reg [31:0] z5681_assgn56814;
    reg [31:0] z5681_assgn56815;
    reg [31:0] z5681_assgn56816;
    reg [31:0] z5681_assgn56817;
    reg [31:0] z5681_assgn56818;
    reg [31:0] z1977_assgn1977;
    wire [31:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p0_0_G16_mul1_G256_inv0;
    wire [31:0] p1_0_G16_mul1_G256_inv0;
    wire [31:0] p0_G16_mul1_G256_inv0;
    wire [31:0] p1_G16_mul1_G256_inv0;
    wire [31:0] z5693_assgn5693;
    reg [31:0] z5693_assgn56930;
    reg [31:0] z5693_assgn56931;
    reg [31:0] z5693_assgn56932;
    reg [31:0] z5693_assgn56933;
    reg [31:0] z5693_assgn56934;
    reg [31:0] z1987_assgn1987;
    wire [31:0] r00_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5697_assgn5697;
    reg [31:0] z5697_assgn56970;
    reg [31:0] z5697_assgn56971;
    reg [31:0] z5697_assgn56972;
    reg [31:0] z5697_assgn56973;
    reg [31:0] z5697_assgn56974;
    reg [31:0] z1989_assgn1989;
    wire [31:0] r10_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5701_assgn5701;
    reg [31:0] z5701_assgn57010;
    reg [31:0] z5701_assgn57011;
    reg [31:0] z5701_assgn57012;
    reg [31:0] z5701_assgn57013;
    reg [31:0] z5701_assgn57014;
    reg [31:0] z1991_assgn1991;
    wire [31:0] r20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5705_assgn5705;
    reg [31:0] z5705_assgn57050;
    reg [31:0] z5705_assgn57051;
    reg [31:0] z5705_assgn57052;
    reg [31:0] z5705_assgn57053;
    reg [31:0] z5705_assgn57054;
    reg [31:0] z5705_assgn57055;
    reg [31:0] z5705_assgn57056;
    reg [31:0] z5705_assgn57057;
    reg [31:0] z1993_assgn1993;
    wire [31:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5709_assgn5709;
    reg [31:0] z5709_assgn57090;
    reg [31:0] z5709_assgn57091;
    reg [31:0] z5709_assgn57092;
    reg [31:0] z5709_assgn57093;
    reg [31:0] z5709_assgn57094;
    reg [31:0] z5709_assgn57095;
    reg [31:0] z5709_assgn57096;
    reg [31:0] z5709_assgn57097;
    reg [31:0] z1995_assgn1995;
    wire [31:0] a1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5713_assgn5713;
    reg [31:0] z5713_assgn57130;
    reg [31:0] z5713_assgn57131;
    reg [31:0] z5713_assgn57132;
    reg [31:0] z5713_assgn57133;
    reg [31:0] z5713_assgn57134;
    reg [31:0] z5713_assgn57135;
    reg [31:0] z5713_assgn57136;
    reg [31:0] z5713_assgn57137;
    reg [31:0] z1997_assgn1997;
    wire [31:0] a0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5717_assgn5717;
    reg [31:0] z5717_assgn57170;
    reg [31:0] z5717_assgn57171;
    reg [31:0] z5717_assgn57172;
    reg [31:0] z5717_assgn57173;
    reg [31:0] z5717_assgn57174;
    reg [31:0] z5717_assgn57175;
    reg [31:0] z5717_assgn57176;
    reg [31:0] z5717_assgn57177;
    reg [31:0] z1999_assgn1999;
    wire [31:0] a1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5721_assgn5721;
    reg [31:0] z5721_assgn57210;
    reg [31:0] z5721_assgn57211;
    reg [31:0] z5721_assgn57212;
    reg [31:0] z5721_assgn57213;
    reg [31:0] z5721_assgn57214;
    reg [31:0] z5721_assgn57215;
    reg [31:0] z5721_assgn57216;
    reg [31:0] z5721_assgn57217;
    reg [31:0] z2001_assgn2001;
    wire [31:0] b0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5725_assgn5725;
    reg [31:0] z5725_assgn57250;
    reg [31:0] z5725_assgn57251;
    reg [31:0] z5725_assgn57252;
    reg [31:0] z5725_assgn57253;
    reg [31:0] z5725_assgn57254;
    reg [31:0] z5725_assgn57255;
    reg [31:0] z5725_assgn57256;
    reg [31:0] z5725_assgn57257;
    reg [31:0] z2003_assgn2003;
    wire [31:0] b1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5729_assgn5729;
    reg [31:0] z5729_assgn57290;
    reg [31:0] z5729_assgn57291;
    reg [31:0] z5729_assgn57292;
    reg [31:0] z5729_assgn57293;
    reg [31:0] z5729_assgn57294;
    reg [31:0] z2005_assgn2005;
    wire [31:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5733_assgn5733;
    reg [31:0] z5733_assgn57330;
    reg [31:0] z5733_assgn57331;
    reg [31:0] z5733_assgn57332;
    reg [31:0] z5733_assgn57333;
    reg [31:0] z5733_assgn57334;
    reg [31:0] z2007_assgn2007;
    wire [31:0] c1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5737_assgn5737;
    reg [31:0] z5737_assgn57370;
    reg [31:0] z5737_assgn57371;
    reg [31:0] z5737_assgn57372;
    reg [31:0] z5737_assgn57373;
    reg [31:0] z5737_assgn57374;
    reg [31:0] z2009_assgn2009;
    wire [31:0] c0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5741_assgn5741;
    reg [31:0] z5741_assgn57410;
    reg [31:0] z5741_assgn57411;
    reg [31:0] z5741_assgn57412;
    reg [31:0] z5741_assgn57413;
    reg [31:0] z5741_assgn57414;
    reg [31:0] z2011_assgn2011;
    wire [31:0] c1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5745_assgn5745;
    reg [31:0] z5745_assgn57450;
    reg [31:0] z5745_assgn57451;
    reg [31:0] z5745_assgn57452;
    reg [31:0] z5745_assgn57453;
    reg [31:0] z5745_assgn57454;
    reg [31:0] z2013_assgn2013;
    wire [31:0] d0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5749_assgn5749;
    reg [31:0] z5749_assgn57490;
    reg [31:0] z5749_assgn57491;
    reg [31:0] z5749_assgn57492;
    reg [31:0] z5749_assgn57493;
    reg [31:0] z5749_assgn57494;
    reg [31:0] z2015_assgn2015;
    wire [31:0] d1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] c0_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] d0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] c1_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] d1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5761_assgn5761;
    reg [31:0] z5761_assgn57610;
    reg [31:0] z5761_assgn57611;
    reg [31:0] z5761_assgn57612;
    reg [31:0] z5761_assgn57613;
    reg [31:0] z5761_assgn57614;
    reg [31:0] z5761_assgn57615;
    reg [31:0] z2025_assgn2025;
    wire [31:0] r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5769_assgn5769;
    reg [31:0] z5769_assgn57690;
    reg [31:0] z2031_assgn2031;
    wire [31:0] u0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5773_assgn5773;
    reg [31:0] z5773_assgn57730;
    reg [31:0] z2033_assgn2033;
    wire [31:0] u1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] cxord_0_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] cxord_1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5781_assgn5781;
    reg [31:0] z5781_assgn57810;
    reg [31:0] z2039_assgn2039;
    wire [31:0] p0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] e0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5791_assgn5791;
    reg [31:0] z5791_assgn57910;
    reg [31:0] z2047_assgn2047;
    wire [31:0] p2_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] e1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5801_assgn5801;
    reg [31:0] z5801_assgn58010;
    reg [31:0] z5801_assgn58011;
    reg [31:0] z5801_assgn58012;
    reg [31:0] z5801_assgn58013;
    reg [31:0] z5801_assgn58014;
    reg [31:0] z5801_assgn58015;
    reg [31:0] z2055_assgn2055;
    wire [31:0] r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5809_assgn5809;
    reg [31:0] z5809_assgn58090;
    reg [31:0] z2061_assgn2061;
    wire [31:0] u0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5813_assgn5813;
    reg [31:0] z5813_assgn58130;
    reg [31:0] z2063_assgn2063;
    wire [31:0] u1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5817_assgn5817;
    reg [31:0] z5817_assgn58170;
    reg [31:0] z2066_assgn2066;
    reg [31:0] r0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5821_assgn5821;
    reg [31:0] z5821_assgn58210;
    reg [31:0] z2068_assgn2068;
    wire [31:0] v1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5825_assgn5825;
    reg [31:0] z5825_assgn58250;
    reg [31:0] z5825_assgn58251;
    reg [31:0] z2069_assgn2069;
    wire [31:0] p0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5835_assgn5835;
    reg [31:0] z5835_assgn58350;
    reg [31:0] z5835_assgn58351;
    reg [31:0] z2077_assgn2077;
    wire [31:0] p2_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5849_assgn5849;
    reg [31:0] z5849_assgn58490;
    reg [31:0] z5849_assgn58491;
    reg [31:0] z5849_assgn58492;
    reg [31:0] z5849_assgn58493;
    reg [31:0] z5849_assgn58494;
    reg [31:0] z5849_assgn58495;
    reg [31:0] z2089_assgn2089;
    wire [31:0] r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5857_assgn5857;
    reg [31:0] z5857_assgn58570;
    reg [31:0] z2095_assgn2095;
    wire [31:0] u0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5861_assgn5861;
    reg [31:0] z5861_assgn58610;
    reg [31:0] z2097_assgn2097;
    wire [31:0] u1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5865_assgn5865;
    reg [31:0] z5865_assgn58650;
    reg [31:0] z2100_assgn2100;
    reg [31:0] r0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5869_assgn5869;
    reg [31:0] z5869_assgn58690;
    reg [31:0] z2102_assgn2102;
    wire [31:0] v1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5873_assgn5873;
    reg [31:0] z5873_assgn58730;
    reg [31:0] z5873_assgn58731;
    reg [31:0] z2103_assgn2103;
    wire [31:0] p0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5883_assgn5883;
    reg [31:0] z5883_assgn58830;
    reg [31:0] z5883_assgn58831;
    reg [31:0] z2111_assgn2111;
    wire [31:0] p2_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5897_assgn5897;
    reg [31:0] z5897_assgn58970;
    reg [31:0] z5897_assgn58971;
    reg [31:0] z5897_assgn58972;
    reg [31:0] z5897_assgn58973;
    reg [31:0] z5897_assgn58974;
    reg [31:0] z5897_assgn58975;
    reg [31:0] z5897_assgn58976;
    reg [31:0] z5897_assgn58977;
    reg [31:0] z5897_assgn58978;
    reg [31:0] z2123_assgn2123;
    wire [31:0] p1ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z5901_assgn5901;
    reg [31:0] z5901_assgn59010;
    reg [31:0] z5901_assgn59011;
    reg [31:0] z5901_assgn59012;
    reg [31:0] z5901_assgn59013;
    reg [31:0] z5901_assgn59014;
    reg [31:0] z5901_assgn59015;
    reg [31:0] z5901_assgn59016;
    reg [31:0] z5901_assgn59017;
    reg [31:0] z5901_assgn59018;
    reg [31:0] z2125_assgn2125;
    wire [31:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q0_0_G16_mul1_G256_inv0;
    wire [31:0] q1_0_G16_mul1_G256_inv0;
    wire [31:0] q0_G16_mul1_G256_inv0;
    wire [31:0] q1_G16_mul1_G256_inv0;
    wire [31:0] z5913_assgn5913;
    reg [31:0] z5913_assgn59130;
    reg [31:0] z5913_assgn59131;
    reg [31:0] z5913_assgn59132;
    reg [31:0] z5913_assgn59133;
    reg [31:0] z5913_assgn59134;
    reg [31:0] z5913_assgn59135;
    reg [31:0] z5913_assgn59136;
    reg [31:0] z5913_assgn59137;
    reg [31:0] z5913_assgn59138;
    reg [31:0] z2135_assgn2135;
    wire [31:0] p0ls2_G16_mul1_G256_inv0;
    wire [31:0] z5917_assgn5917;
    reg [31:0] z5917_assgn59170;
    reg [31:0] z5917_assgn59171;
    reg [31:0] z5917_assgn59172;
    reg [31:0] z5917_assgn59173;
    reg [31:0] z5917_assgn59174;
    reg [31:0] z5917_assgn59175;
    reg [31:0] z5917_assgn59176;
    reg [31:0] z5917_assgn59177;
    reg [31:0] z5917_assgn59178;
    reg [31:0] z2137_assgn2137;
    wire [31:0] p1ls2_G16_mul1_G256_inv0;
    wire [31:0] p0_G256_inv0;
    wire [31:0] p1_G256_inv0;
    wire [31:0] z5925_assgn5925;
    reg [31:0] z5925_assgn59250;
    reg [31:0] z5925_assgn59251;
    reg [31:0] z5925_assgn59252;
    reg [31:0] z5925_assgn59253;
    reg [31:0] z5925_assgn59254;
    reg [31:0] z2143_assgn2143;
    wire [31:0] r00_G16_mul2_G256_inv0;
    wire [31:0] z5929_assgn5929;
    reg [31:0] z5929_assgn59290;
    reg [31:0] z5929_assgn59291;
    reg [31:0] z5929_assgn59292;
    reg [31:0] z5929_assgn59293;
    reg [31:0] z5929_assgn59294;
    reg [31:0] z2145_assgn2145;
    wire [31:0] r10_G16_mul2_G256_inv0;
    wire [31:0] z5933_assgn5933;
    reg [31:0] z5933_assgn59330;
    reg [31:0] z5933_assgn59331;
    reg [31:0] z5933_assgn59332;
    reg [31:0] z5933_assgn59333;
    reg [31:0] z5933_assgn59334;
    reg [31:0] z2147_assgn2147;
    wire [31:0] r20_G16_mul2_G256_inv0;
    wire [31:0] z5937_assgn5937;
    reg [31:0] z5937_assgn59370;
    reg [31:0] z5937_assgn59371;
    reg [31:0] z5937_assgn59372;
    reg [31:0] z5937_assgn59373;
    reg [31:0] z5937_assgn59374;
    reg [31:0] z2149_assgn2149;
    wire [31:0] r30_G16_mul2_G256_inv0;
    wire [31:0] z5941_assgn5941;
    reg [31:0] z5941_assgn59410;
    reg [31:0] z5941_assgn59411;
    reg [31:0] z5941_assgn59412;
    reg [31:0] z5941_assgn59413;
    reg [31:0] z5941_assgn59414;
    reg [31:0] z2151_assgn2151;
    wire [31:0] r40_G16_mul2_G256_inv0;
    wire [31:0] z5945_assgn5945;
    reg [31:0] z5945_assgn59450;
    reg [31:0] z5945_assgn59451;
    reg [31:0] z5945_assgn59452;
    reg [31:0] z5945_assgn59453;
    reg [31:0] z5945_assgn59454;
    reg [31:0] z2153_assgn2153;
    wire [31:0] r50_G16_mul2_G256_inv0;
    wire [31:0] z5949_assgn5949;
    reg [31:0] z5949_assgn59490;
    reg [31:0] z5949_assgn59491;
    reg [31:0] z5949_assgn59492;
    reg [31:0] z5949_assgn59493;
    reg [31:0] z5949_assgn59494;
    reg [31:0] z2155_assgn2155;
    wire [31:0] r60_G16_mul2_G256_inv0;
    wire [31:0] z5953_assgn5953;
    reg [31:0] z5953_assgn59530;
    reg [31:0] z5953_assgn59531;
    reg [31:0] z5953_assgn59532;
    reg [31:0] z5953_assgn59533;
    reg [31:0] z5953_assgn59534;
    reg [31:0] z2157_assgn2157;
    wire [31:0] r70_G16_mul2_G256_inv0;
    wire [31:0] z5957_assgn5957;
    reg [31:0] z5957_assgn59570;
    reg [31:0] z5957_assgn59571;
    reg [31:0] z5957_assgn59572;
    reg [31:0] z5957_assgn59573;
    reg [31:0] z5957_assgn59574;
    reg [31:0] z2159_assgn2159;
    wire [31:0] r80_G16_mul2_G256_inv0;
    wire [31:0] z5961_assgn5961;
    reg [31:0] z5961_assgn59610;
    reg [31:0] z5961_assgn59611;
    reg [31:0] z5961_assgn59612;
    reg [31:0] z5961_assgn59613;
    reg [31:0] z5961_assgn59614;
    reg [31:0] z5961_assgn59615;
    reg [31:0] z5961_assgn59616;
    reg [31:0] z5961_assgn59617;
    reg [31:0] z2161_assgn2161;
    wire [31:0] a0_0_G16_mul2_G256_inv0;
    wire [31:0] z5965_assgn5965;
    reg [31:0] z5965_assgn59650;
    reg [31:0] z5965_assgn59651;
    reg [31:0] z5965_assgn59652;
    reg [31:0] z5965_assgn59653;
    reg [31:0] z5965_assgn59654;
    reg [31:0] z5965_assgn59655;
    reg [31:0] z5965_assgn59656;
    reg [31:0] z5965_assgn59657;
    reg [31:0] z2163_assgn2163;
    wire [31:0] a1_0_G16_mul2_G256_inv0;
    wire [31:0] z5969_assgn5969;
    reg [31:0] z5969_assgn59690;
    reg [31:0] z5969_assgn59691;
    reg [31:0] z5969_assgn59692;
    reg [31:0] z5969_assgn59693;
    reg [31:0] z5969_assgn59694;
    reg [31:0] z5969_assgn59695;
    reg [31:0] z5969_assgn59696;
    reg [31:0] z5969_assgn59697;
    reg [31:0] z2165_assgn2165;
    wire [31:0] a0_G16_mul2_G256_inv0;
    wire [31:0] z5973_assgn5973;
    reg [31:0] z5973_assgn59730;
    reg [31:0] z5973_assgn59731;
    reg [31:0] z5973_assgn59732;
    reg [31:0] z5973_assgn59733;
    reg [31:0] z5973_assgn59734;
    reg [31:0] z5973_assgn59735;
    reg [31:0] z5973_assgn59736;
    reg [31:0] z5973_assgn59737;
    reg [31:0] z2167_assgn2167;
    wire [31:0] a1_G16_mul2_G256_inv0;
    wire [31:0] z5977_assgn5977;
    reg [31:0] z5977_assgn59770;
    reg [31:0] z5977_assgn59771;
    reg [31:0] z5977_assgn59772;
    reg [31:0] z5977_assgn59773;
    reg [31:0] z5977_assgn59774;
    reg [31:0] z5977_assgn59775;
    reg [31:0] z5977_assgn59776;
    reg [31:0] z5977_assgn59777;
    reg [31:0] z2169_assgn2169;
    wire [31:0] b0_G16_mul2_G256_inv0;
    wire [31:0] z5981_assgn5981;
    reg [31:0] z5981_assgn59810;
    reg [31:0] z5981_assgn59811;
    reg [31:0] z5981_assgn59812;
    reg [31:0] z5981_assgn59813;
    reg [31:0] z5981_assgn59814;
    reg [31:0] z5981_assgn59815;
    reg [31:0] z5981_assgn59816;
    reg [31:0] z5981_assgn59817;
    reg [31:0] z2171_assgn2171;
    wire [31:0] b1_G16_mul2_G256_inv0;
    wire [31:0] z5985_assgn5985;
    reg [31:0] z5985_assgn59850;
    reg [31:0] z5985_assgn59851;
    reg [31:0] z5985_assgn59852;
    reg [31:0] z5985_assgn59853;
    reg [31:0] z5985_assgn59854;
    reg [31:0] z2173_assgn2173;
    wire [31:0] z5987_assgn5987;
    reg [31:0] z5987_assgn59870;
    reg [31:0] z5987_assgn59871;
    reg [31:0] z2174_assgn2174;
    wire [31:0] c0_0_G16_mul2_G256_inv0;
    wire [31:0] z5991_assgn5991;
    reg [31:0] z5991_assgn59910;
    reg [31:0] z5991_assgn59911;
    reg [31:0] z5991_assgn59912;
    reg [31:0] z5991_assgn59913;
    reg [31:0] z5991_assgn59914;
    reg [31:0] z2175_assgn2175;
    wire [31:0] z5993_assgn5993;
    reg [31:0] z5993_assgn59930;
    reg [31:0] z5993_assgn59931;
    reg [31:0] z2176_assgn2176;
    wire [31:0] c1_0_G16_mul2_G256_inv0;
    wire [31:0] z5997_assgn5997;
    reg [31:0] z5997_assgn59970;
    reg [31:0] z5997_assgn59971;
    reg [31:0] z5997_assgn59972;
    reg [31:0] z5997_assgn59973;
    reg [31:0] z5997_assgn59974;
    reg [31:0] z2177_assgn2177;
    wire [31:0] c0_G16_mul2_G256_inv0;
    wire [31:0] z6001_assgn6001;
    reg [31:0] z6001_assgn60010;
    reg [31:0] z6001_assgn60011;
    reg [31:0] z6001_assgn60012;
    reg [31:0] z6001_assgn60013;
    reg [31:0] z6001_assgn60014;
    reg [31:0] z2179_assgn2179;
    wire [31:0] c1_G16_mul2_G256_inv0;
    wire [31:0] z6005_assgn6005;
    reg [31:0] z6005_assgn60050;
    reg [31:0] z6005_assgn60051;
    reg [31:0] z6005_assgn60052;
    reg [31:0] z6005_assgn60053;
    reg [31:0] z6005_assgn60054;
    reg [31:0] z2181_assgn2181;
    wire [31:0] z6007_assgn6007;
    reg [31:0] z6007_assgn60070;
    reg [31:0] z6007_assgn60071;
    reg [31:0] z2182_assgn2182;
    wire [31:0] d0_G16_mul2_G256_inv0;
    wire [31:0] z6011_assgn6011;
    reg [31:0] z6011_assgn60110;
    reg [31:0] z6011_assgn60111;
    reg [31:0] z6011_assgn60112;
    reg [31:0] z6011_assgn60113;
    reg [31:0] z6011_assgn60114;
    reg [31:0] z2183_assgn2183;
    wire [31:0] z6013_assgn6013;
    reg [31:0] z6013_assgn60130;
    reg [31:0] z6013_assgn60131;
    reg [31:0] z2184_assgn2184;
    wire [31:0] d1_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G16_mul2_G256_inv0;
    wire [31:0] cxord_0_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G16_mul2_G256_inv0;
    wire [31:0] cxord_1_G16_mul2_G256_inv0;
    wire [31:0] z6025_assgn6025;
    reg [31:0] z6025_assgn60250;
    reg [31:0] z6025_assgn60251;
    reg [31:0] z6025_assgn60252;
    reg [31:0] z6025_assgn60253;
    reg [31:0] z6025_assgn60254;
    reg [31:0] z2193_assgn2193;
    wire [31:0] r00_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6029_assgn6029;
    reg [31:0] z6029_assgn60290;
    reg [31:0] z6029_assgn60291;
    reg [31:0] z6029_assgn60292;
    reg [31:0] z6029_assgn60293;
    reg [31:0] z6029_assgn60294;
    reg [31:0] z2195_assgn2195;
    wire [31:0] r10_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6033_assgn6033;
    reg [31:0] z6033_assgn60330;
    reg [31:0] z6033_assgn60331;
    reg [31:0] z6033_assgn60332;
    reg [31:0] z6033_assgn60333;
    reg [31:0] z6033_assgn60334;
    reg [31:0] z2197_assgn2197;
    wire [31:0] r20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6037_assgn6037;
    reg [31:0] z6037_assgn60370;
    reg [31:0] z6037_assgn60371;
    reg [31:0] z6037_assgn60372;
    reg [31:0] z6037_assgn60373;
    reg [31:0] z6037_assgn60374;
    reg [31:0] z6037_assgn60375;
    reg [31:0] z6037_assgn60376;
    reg [31:0] z6037_assgn60377;
    reg [31:0] z2199_assgn2199;
    wire [31:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6041_assgn6041;
    reg [31:0] z6041_assgn60410;
    reg [31:0] z6041_assgn60411;
    reg [31:0] z6041_assgn60412;
    reg [31:0] z6041_assgn60413;
    reg [31:0] z6041_assgn60414;
    reg [31:0] z6041_assgn60415;
    reg [31:0] z6041_assgn60416;
    reg [31:0] z6041_assgn60417;
    reg [31:0] z2201_assgn2201;
    wire [31:0] a1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6045_assgn6045;
    reg [31:0] z6045_assgn60450;
    reg [31:0] z6045_assgn60451;
    reg [31:0] z6045_assgn60452;
    reg [31:0] z6045_assgn60453;
    reg [31:0] z6045_assgn60454;
    reg [31:0] z6045_assgn60455;
    reg [31:0] z6045_assgn60456;
    reg [31:0] z6045_assgn60457;
    reg [31:0] z2203_assgn2203;
    wire [31:0] a0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6049_assgn6049;
    reg [31:0] z6049_assgn60490;
    reg [31:0] z6049_assgn60491;
    reg [31:0] z6049_assgn60492;
    reg [31:0] z6049_assgn60493;
    reg [31:0] z6049_assgn60494;
    reg [31:0] z6049_assgn60495;
    reg [31:0] z6049_assgn60496;
    reg [31:0] z6049_assgn60497;
    reg [31:0] z2205_assgn2205;
    wire [31:0] a1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6053_assgn6053;
    reg [31:0] z6053_assgn60530;
    reg [31:0] z6053_assgn60531;
    reg [31:0] z6053_assgn60532;
    reg [31:0] z6053_assgn60533;
    reg [31:0] z6053_assgn60534;
    reg [31:0] z6053_assgn60535;
    reg [31:0] z6053_assgn60536;
    reg [31:0] z6053_assgn60537;
    reg [31:0] z2207_assgn2207;
    wire [31:0] b0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6057_assgn6057;
    reg [31:0] z6057_assgn60570;
    reg [31:0] z6057_assgn60571;
    reg [31:0] z6057_assgn60572;
    reg [31:0] z6057_assgn60573;
    reg [31:0] z6057_assgn60574;
    reg [31:0] z6057_assgn60575;
    reg [31:0] z6057_assgn60576;
    reg [31:0] z6057_assgn60577;
    reg [31:0] z2209_assgn2209;
    wire [31:0] b1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6061_assgn6061;
    reg [31:0] z6061_assgn60610;
    reg [31:0] z6061_assgn60611;
    reg [31:0] z6061_assgn60612;
    reg [31:0] z6061_assgn60613;
    reg [31:0] z6061_assgn60614;
    reg [31:0] z2211_assgn2211;
    wire [31:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6065_assgn6065;
    reg [31:0] z6065_assgn60650;
    reg [31:0] z6065_assgn60651;
    reg [31:0] z6065_assgn60652;
    reg [31:0] z6065_assgn60653;
    reg [31:0] z6065_assgn60654;
    reg [31:0] z2213_assgn2213;
    wire [31:0] c1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6069_assgn6069;
    reg [31:0] z6069_assgn60690;
    reg [31:0] z6069_assgn60691;
    reg [31:0] z6069_assgn60692;
    reg [31:0] z6069_assgn60693;
    reg [31:0] z6069_assgn60694;
    reg [31:0] z2215_assgn2215;
    wire [31:0] c0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6073_assgn6073;
    reg [31:0] z6073_assgn60730;
    reg [31:0] z6073_assgn60731;
    reg [31:0] z6073_assgn60732;
    reg [31:0] z6073_assgn60733;
    reg [31:0] z6073_assgn60734;
    reg [31:0] z2217_assgn2217;
    wire [31:0] c1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6077_assgn6077;
    reg [31:0] z6077_assgn60770;
    reg [31:0] z6077_assgn60771;
    reg [31:0] z6077_assgn60772;
    reg [31:0] z6077_assgn60773;
    reg [31:0] z6077_assgn60774;
    reg [31:0] z2219_assgn2219;
    wire [31:0] d0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6081_assgn6081;
    reg [31:0] z6081_assgn60810;
    reg [31:0] z6081_assgn60811;
    reg [31:0] z6081_assgn60812;
    reg [31:0] z6081_assgn60813;
    reg [31:0] z6081_assgn60814;
    reg [31:0] z2221_assgn2221;
    wire [31:0] d1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] c0_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] d0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] c1_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] d1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6093_assgn6093;
    reg [31:0] z6093_assgn60930;
    reg [31:0] z6093_assgn60931;
    reg [31:0] z6093_assgn60932;
    reg [31:0] z6093_assgn60933;
    reg [31:0] z6093_assgn60934;
    reg [31:0] z6093_assgn60935;
    reg [31:0] z2231_assgn2231;
    wire [31:0] r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6101_assgn6101;
    reg [31:0] z6101_assgn61010;
    reg [31:0] z2237_assgn2237;
    wire [31:0] u0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6105_assgn6105;
    reg [31:0] z6105_assgn61050;
    reg [31:0] z2239_assgn2239;
    wire [31:0] u1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] cxord_0_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] cxord_1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6113_assgn6113;
    reg [31:0] z6113_assgn61130;
    reg [31:0] z2245_assgn2245;
    wire [31:0] p0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] e0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6123_assgn6123;
    reg [31:0] z6123_assgn61230;
    reg [31:0] z2253_assgn2253;
    wire [31:0] p2_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] e1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6133_assgn6133;
    reg [31:0] z6133_assgn61330;
    reg [31:0] z6133_assgn61331;
    reg [31:0] z6133_assgn61332;
    reg [31:0] z6133_assgn61333;
    reg [31:0] z6133_assgn61334;
    reg [31:0] z6133_assgn61335;
    reg [31:0] z2261_assgn2261;
    wire [31:0] r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6141_assgn6141;
    reg [31:0] z6141_assgn61410;
    reg [31:0] z2267_assgn2267;
    wire [31:0] u0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6145_assgn6145;
    reg [31:0] z6145_assgn61450;
    reg [31:0] z2269_assgn2269;
    wire [31:0] u1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6149_assgn6149;
    reg [31:0] z6149_assgn61490;
    reg [31:0] z2272_assgn2272;
    reg [31:0] r0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6153_assgn6153;
    reg [31:0] z6153_assgn61530;
    reg [31:0] z2274_assgn2274;
    wire [31:0] v1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6157_assgn6157;
    reg [31:0] z6157_assgn61570;
    reg [31:0] z6157_assgn61571;
    reg [31:0] z2275_assgn2275;
    wire [31:0] p0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6167_assgn6167;
    reg [31:0] z6167_assgn61670;
    reg [31:0] z6167_assgn61671;
    reg [31:0] z2283_assgn2283;
    wire [31:0] p2_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6181_assgn6181;
    reg [31:0] z6181_assgn61810;
    reg [31:0] z6181_assgn61811;
    reg [31:0] z6181_assgn61812;
    reg [31:0] z6181_assgn61813;
    reg [31:0] z6181_assgn61814;
    reg [31:0] z6181_assgn61815;
    reg [31:0] z2295_assgn2295;
    wire [31:0] r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6189_assgn6189;
    reg [31:0] z6189_assgn61890;
    reg [31:0] z2301_assgn2301;
    wire [31:0] u0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6193_assgn6193;
    reg [31:0] z6193_assgn61930;
    reg [31:0] z2303_assgn2303;
    wire [31:0] u1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6197_assgn6197;
    reg [31:0] z6197_assgn61970;
    reg [31:0] z2306_assgn2306;
    reg [31:0] r0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6201_assgn6201;
    reg [31:0] z6201_assgn62010;
    reg [31:0] z2308_assgn2308;
    wire [31:0] v1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6205_assgn6205;
    reg [31:0] z6205_assgn62050;
    reg [31:0] z6205_assgn62051;
    reg [31:0] z2309_assgn2309;
    wire [31:0] p0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6215_assgn6215;
    reg [31:0] z6215_assgn62150;
    reg [31:0] z6215_assgn62151;
    reg [31:0] z2317_assgn2317;
    wire [31:0] p2_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6229_assgn6229;
    reg [31:0] z6229_assgn62290;
    reg [31:0] z6229_assgn62291;
    reg [31:0] z6229_assgn62292;
    reg [31:0] z6229_assgn62293;
    reg [31:0] z6229_assgn62294;
    reg [31:0] z6229_assgn62295;
    reg [31:0] z6229_assgn62296;
    reg [31:0] z6229_assgn62297;
    reg [31:0] z6229_assgn62298;
    reg [31:0] z2329_assgn2329;
    wire [31:0] p1ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6233_assgn6233;
    reg [31:0] z6233_assgn62330;
    reg [31:0] z6233_assgn62331;
    reg [31:0] z6233_assgn62332;
    reg [31:0] z6233_assgn62333;
    reg [31:0] z6233_assgn62334;
    reg [31:0] z6233_assgn62335;
    reg [31:0] z6233_assgn62336;
    reg [31:0] z6233_assgn62337;
    reg [31:0] z6233_assgn62338;
    reg [31:0] z2331_assgn2331;
    wire [31:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] e0_G16_mul2_G256_inv0;
    wire [31:0] e1_G16_mul2_G256_inv0;
    wire [31:0] z6241_assgn6241;
    reg [31:0] z6241_assgn62410;
    reg [31:0] z6241_assgn62411;
    reg [31:0] z6241_assgn62412;
    reg [31:0] z6241_assgn62413;
    reg [31:0] z6241_assgn62414;
    reg [31:0] z6241_assgn62415;
    reg [31:0] z6241_assgn62416;
    reg [31:0] z6241_assgn62417;
    reg [31:0] z6241_assgn62418;
    reg [31:0] z2337_assgn2337;
    wire [31:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6245_assgn6245;
    reg [31:0] z6245_assgn62450;
    reg [31:0] z6245_assgn62451;
    reg [31:0] z6245_assgn62452;
    reg [31:0] z6245_assgn62453;
    reg [31:0] z6245_assgn62454;
    reg [31:0] z6245_assgn62455;
    reg [31:0] z6245_assgn62456;
    reg [31:0] z6245_assgn62457;
    reg [31:0] z6245_assgn62458;
    reg [31:0] z2339_assgn2339;
    wire [31:0] a1_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6249_assgn6249;
    reg [31:0] z6249_assgn62490;
    reg [31:0] z6249_assgn62491;
    reg [31:0] z6249_assgn62492;
    reg [31:0] z6249_assgn62493;
    reg [31:0] z6249_assgn62494;
    reg [31:0] z6249_assgn62495;
    reg [31:0] z6249_assgn62496;
    reg [31:0] z6249_assgn62497;
    reg [31:0] z6249_assgn62498;
    reg [31:0] z2341_assgn2341;
    wire [31:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6253_assgn6253;
    reg [31:0] z6253_assgn62530;
    reg [31:0] z6253_assgn62531;
    reg [31:0] z6253_assgn62532;
    reg [31:0] z6253_assgn62533;
    reg [31:0] z6253_assgn62534;
    reg [31:0] z6253_assgn62535;
    reg [31:0] z6253_assgn62536;
    reg [31:0] z6253_assgn62537;
    reg [31:0] z6253_assgn62538;
    reg [31:0] z2343_assgn2343;
    wire [31:0] a1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6257_assgn6257;
    reg [31:0] z6257_assgn62570;
    reg [31:0] z6257_assgn62571;
    reg [31:0] z6257_assgn62572;
    reg [31:0] z6257_assgn62573;
    reg [31:0] z6257_assgn62574;
    reg [31:0] z6257_assgn62575;
    reg [31:0] z6257_assgn62576;
    reg [31:0] z6257_assgn62577;
    reg [31:0] z6257_assgn62578;
    reg [31:0] z2345_assgn2345;
    wire [31:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6261_assgn6261;
    reg [31:0] z6261_assgn62610;
    reg [31:0] z6261_assgn62611;
    reg [31:0] z6261_assgn62612;
    reg [31:0] z6261_assgn62613;
    reg [31:0] z6261_assgn62614;
    reg [31:0] z6261_assgn62615;
    reg [31:0] z6261_assgn62616;
    reg [31:0] z6261_assgn62617;
    reg [31:0] z6261_assgn62618;
    reg [31:0] z2347_assgn2347;
    wire [31:0] b1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6273_assgn6273;
    reg [31:0] z6273_assgn62730;
    reg [31:0] z6273_assgn62731;
    reg [31:0] z6273_assgn62732;
    reg [31:0] z6273_assgn62733;
    reg [31:0] z6273_assgn62734;
    reg [31:0] z6273_assgn62735;
    reg [31:0] z6273_assgn62736;
    reg [31:0] z6273_assgn62737;
    reg [31:0] z6273_assgn62738;
    reg [31:0] z2357_assgn2357;
    wire [31:0] p1ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z6277_assgn6277;
    reg [31:0] z6277_assgn62770;
    reg [31:0] z6277_assgn62771;
    reg [31:0] z6277_assgn62772;
    reg [31:0] z6277_assgn62773;
    reg [31:0] z6277_assgn62774;
    reg [31:0] z6277_assgn62775;
    reg [31:0] z6277_assgn62776;
    reg [31:0] z6277_assgn62777;
    reg [31:0] z6277_assgn62778;
    reg [31:0] z2359_assgn2359;
    wire [31:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] e01_G16_mul2_G256_inv0;
    wire [31:0] e11_G16_mul2_G256_inv0;
    wire [31:0] z6285_assgn6285;
    reg [31:0] z6285_assgn62850;
    reg [31:0] z6285_assgn62851;
    reg [31:0] z6285_assgn62852;
    reg [31:0] z6285_assgn62853;
    reg [31:0] z6285_assgn62854;
    reg [31:0] z2365_assgn2365;
    wire [31:0] r00_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6289_assgn6289;
    reg [31:0] z6289_assgn62890;
    reg [31:0] z6289_assgn62891;
    reg [31:0] z6289_assgn62892;
    reg [31:0] z6289_assgn62893;
    reg [31:0] z6289_assgn62894;
    reg [31:0] z2367_assgn2367;
    wire [31:0] r10_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6293_assgn6293;
    reg [31:0] z6293_assgn62930;
    reg [31:0] z6293_assgn62931;
    reg [31:0] z6293_assgn62932;
    reg [31:0] z6293_assgn62933;
    reg [31:0] z6293_assgn62934;
    reg [31:0] z2369_assgn2369;
    wire [31:0] r20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6297_assgn6297;
    reg [31:0] z6297_assgn62970;
    reg [31:0] z6297_assgn62971;
    reg [31:0] z6297_assgn62972;
    reg [31:0] z6297_assgn62973;
    reg [31:0] z6297_assgn62974;
    reg [31:0] z6297_assgn62975;
    reg [31:0] z6297_assgn62976;
    reg [31:0] z6297_assgn62977;
    reg [31:0] z2371_assgn2371;
    wire [31:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6301_assgn6301;
    reg [31:0] z6301_assgn63010;
    reg [31:0] z6301_assgn63011;
    reg [31:0] z6301_assgn63012;
    reg [31:0] z6301_assgn63013;
    reg [31:0] z6301_assgn63014;
    reg [31:0] z6301_assgn63015;
    reg [31:0] z6301_assgn63016;
    reg [31:0] z6301_assgn63017;
    reg [31:0] z2373_assgn2373;
    wire [31:0] a1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6305_assgn6305;
    reg [31:0] z6305_assgn63050;
    reg [31:0] z6305_assgn63051;
    reg [31:0] z6305_assgn63052;
    reg [31:0] z6305_assgn63053;
    reg [31:0] z6305_assgn63054;
    reg [31:0] z6305_assgn63055;
    reg [31:0] z6305_assgn63056;
    reg [31:0] z6305_assgn63057;
    reg [31:0] z2375_assgn2375;
    wire [31:0] a0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6309_assgn6309;
    reg [31:0] z6309_assgn63090;
    reg [31:0] z6309_assgn63091;
    reg [31:0] z6309_assgn63092;
    reg [31:0] z6309_assgn63093;
    reg [31:0] z6309_assgn63094;
    reg [31:0] z6309_assgn63095;
    reg [31:0] z6309_assgn63096;
    reg [31:0] z6309_assgn63097;
    reg [31:0] z2377_assgn2377;
    wire [31:0] a1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6313_assgn6313;
    reg [31:0] z6313_assgn63130;
    reg [31:0] z6313_assgn63131;
    reg [31:0] z6313_assgn63132;
    reg [31:0] z6313_assgn63133;
    reg [31:0] z6313_assgn63134;
    reg [31:0] z6313_assgn63135;
    reg [31:0] z6313_assgn63136;
    reg [31:0] z6313_assgn63137;
    reg [31:0] z2379_assgn2379;
    wire [31:0] b0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6317_assgn6317;
    reg [31:0] z6317_assgn63170;
    reg [31:0] z6317_assgn63171;
    reg [31:0] z6317_assgn63172;
    reg [31:0] z6317_assgn63173;
    reg [31:0] z6317_assgn63174;
    reg [31:0] z6317_assgn63175;
    reg [31:0] z6317_assgn63176;
    reg [31:0] z6317_assgn63177;
    reg [31:0] z2381_assgn2381;
    wire [31:0] b1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6321_assgn6321;
    reg [31:0] z6321_assgn63210;
    reg [31:0] z6321_assgn63211;
    reg [31:0] z6321_assgn63212;
    reg [31:0] z6321_assgn63213;
    reg [31:0] z6321_assgn63214;
    reg [31:0] z2383_assgn2383;
    wire [31:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6325_assgn6325;
    reg [31:0] z6325_assgn63250;
    reg [31:0] z6325_assgn63251;
    reg [31:0] z6325_assgn63252;
    reg [31:0] z6325_assgn63253;
    reg [31:0] z6325_assgn63254;
    reg [31:0] z2385_assgn2385;
    wire [31:0] c1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6329_assgn6329;
    reg [31:0] z6329_assgn63290;
    reg [31:0] z6329_assgn63291;
    reg [31:0] z6329_assgn63292;
    reg [31:0] z6329_assgn63293;
    reg [31:0] z6329_assgn63294;
    reg [31:0] z2387_assgn2387;
    wire [31:0] c0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6333_assgn6333;
    reg [31:0] z6333_assgn63330;
    reg [31:0] z6333_assgn63331;
    reg [31:0] z6333_assgn63332;
    reg [31:0] z6333_assgn63333;
    reg [31:0] z6333_assgn63334;
    reg [31:0] z2389_assgn2389;
    wire [31:0] c1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6337_assgn6337;
    reg [31:0] z6337_assgn63370;
    reg [31:0] z6337_assgn63371;
    reg [31:0] z6337_assgn63372;
    reg [31:0] z6337_assgn63373;
    reg [31:0] z6337_assgn63374;
    reg [31:0] z2391_assgn2391;
    wire [31:0] d0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6341_assgn6341;
    reg [31:0] z6341_assgn63410;
    reg [31:0] z6341_assgn63411;
    reg [31:0] z6341_assgn63412;
    reg [31:0] z6341_assgn63413;
    reg [31:0] z6341_assgn63414;
    reg [31:0] z2393_assgn2393;
    wire [31:0] d1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] c0_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] d0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] c1_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] d1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6353_assgn6353;
    reg [31:0] z6353_assgn63530;
    reg [31:0] z6353_assgn63531;
    reg [31:0] z6353_assgn63532;
    reg [31:0] z6353_assgn63533;
    reg [31:0] z6353_assgn63534;
    reg [31:0] z6353_assgn63535;
    reg [31:0] z2403_assgn2403;
    wire [31:0] r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6361_assgn6361;
    reg [31:0] z6361_assgn63610;
    reg [31:0] z2409_assgn2409;
    wire [31:0] u0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6365_assgn6365;
    reg [31:0] z6365_assgn63650;
    reg [31:0] z2411_assgn2411;
    wire [31:0] u1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] cxord_0_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] cxord_1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6373_assgn6373;
    reg [31:0] z6373_assgn63730;
    reg [31:0] z2417_assgn2417;
    wire [31:0] p0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] e0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6383_assgn6383;
    reg [31:0] z6383_assgn63830;
    reg [31:0] z2425_assgn2425;
    wire [31:0] p2_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] e1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6393_assgn6393;
    reg [31:0] z6393_assgn63930;
    reg [31:0] z6393_assgn63931;
    reg [31:0] z6393_assgn63932;
    reg [31:0] z6393_assgn63933;
    reg [31:0] z6393_assgn63934;
    reg [31:0] z6393_assgn63935;
    reg [31:0] z2433_assgn2433;
    wire [31:0] r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6401_assgn6401;
    reg [31:0] z6401_assgn64010;
    reg [31:0] z2439_assgn2439;
    wire [31:0] u0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6405_assgn6405;
    reg [31:0] z6405_assgn64050;
    reg [31:0] z2441_assgn2441;
    wire [31:0] u1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6409_assgn6409;
    reg [31:0] z6409_assgn64090;
    reg [31:0] z2444_assgn2444;
    reg [31:0] r0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6413_assgn6413;
    reg [31:0] z6413_assgn64130;
    reg [31:0] z2446_assgn2446;
    wire [31:0] v1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6417_assgn6417;
    reg [31:0] z6417_assgn64170;
    reg [31:0] z6417_assgn64171;
    reg [31:0] z2447_assgn2447;
    wire [31:0] p0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6427_assgn6427;
    reg [31:0] z6427_assgn64270;
    reg [31:0] z6427_assgn64271;
    reg [31:0] z2455_assgn2455;
    wire [31:0] p2_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6441_assgn6441;
    reg [31:0] z6441_assgn64410;
    reg [31:0] z6441_assgn64411;
    reg [31:0] z6441_assgn64412;
    reg [31:0] z6441_assgn64413;
    reg [31:0] z6441_assgn64414;
    reg [31:0] z6441_assgn64415;
    reg [31:0] z2467_assgn2467;
    wire [31:0] r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6449_assgn6449;
    reg [31:0] z6449_assgn64490;
    reg [31:0] z2473_assgn2473;
    wire [31:0] u0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6453_assgn6453;
    reg [31:0] z6453_assgn64530;
    reg [31:0] z2475_assgn2475;
    wire [31:0] u1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6457_assgn6457;
    reg [31:0] z6457_assgn64570;
    reg [31:0] z2478_assgn2478;
    reg [31:0] r0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6461_assgn6461;
    reg [31:0] z6461_assgn64610;
    reg [31:0] z2480_assgn2480;
    wire [31:0] v1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6465_assgn6465;
    reg [31:0] z6465_assgn64650;
    reg [31:0] z6465_assgn64651;
    reg [31:0] z2481_assgn2481;
    wire [31:0] p0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6475_assgn6475;
    reg [31:0] z6475_assgn64750;
    reg [31:0] z6475_assgn64751;
    reg [31:0] z2489_assgn2489;
    wire [31:0] p2_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6489_assgn6489;
    reg [31:0] z6489_assgn64890;
    reg [31:0] z6489_assgn64891;
    reg [31:0] z6489_assgn64892;
    reg [31:0] z6489_assgn64893;
    reg [31:0] z6489_assgn64894;
    reg [31:0] z6489_assgn64895;
    reg [31:0] z6489_assgn64896;
    reg [31:0] z6489_assgn64897;
    reg [31:0] z6489_assgn64898;
    reg [31:0] z2501_assgn2501;
    wire [31:0] p1ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z6493_assgn6493;
    reg [31:0] z6493_assgn64930;
    reg [31:0] z6493_assgn64931;
    reg [31:0] z6493_assgn64932;
    reg [31:0] z6493_assgn64933;
    reg [31:0] z6493_assgn64934;
    reg [31:0] z6493_assgn64935;
    reg [31:0] z6493_assgn64936;
    reg [31:0] z6493_assgn64937;
    reg [31:0] z6493_assgn64938;
    reg [31:0] z2503_assgn2503;
    wire [31:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p0_0_G16_mul2_G256_inv0;
    wire [31:0] p1_0_G16_mul2_G256_inv0;
    wire [31:0] p0_G16_mul2_G256_inv0;
    wire [31:0] p1_G16_mul2_G256_inv0;
    wire [31:0] z6505_assgn6505;
    reg [31:0] z6505_assgn65050;
    reg [31:0] z6505_assgn65051;
    reg [31:0] z6505_assgn65052;
    reg [31:0] z6505_assgn65053;
    reg [31:0] z6505_assgn65054;
    reg [31:0] z2513_assgn2513;
    wire [31:0] r00_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6509_assgn6509;
    reg [31:0] z6509_assgn65090;
    reg [31:0] z6509_assgn65091;
    reg [31:0] z6509_assgn65092;
    reg [31:0] z6509_assgn65093;
    reg [31:0] z6509_assgn65094;
    reg [31:0] z2515_assgn2515;
    wire [31:0] r10_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6513_assgn6513;
    reg [31:0] z6513_assgn65130;
    reg [31:0] z6513_assgn65131;
    reg [31:0] z6513_assgn65132;
    reg [31:0] z6513_assgn65133;
    reg [31:0] z6513_assgn65134;
    reg [31:0] z2517_assgn2517;
    wire [31:0] r20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6517_assgn6517;
    reg [31:0] z6517_assgn65170;
    reg [31:0] z6517_assgn65171;
    reg [31:0] z6517_assgn65172;
    reg [31:0] z6517_assgn65173;
    reg [31:0] z6517_assgn65174;
    reg [31:0] z6517_assgn65175;
    reg [31:0] z6517_assgn65176;
    reg [31:0] z6517_assgn65177;
    reg [31:0] z2519_assgn2519;
    wire [31:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6521_assgn6521;
    reg [31:0] z6521_assgn65210;
    reg [31:0] z6521_assgn65211;
    reg [31:0] z6521_assgn65212;
    reg [31:0] z6521_assgn65213;
    reg [31:0] z6521_assgn65214;
    reg [31:0] z6521_assgn65215;
    reg [31:0] z6521_assgn65216;
    reg [31:0] z6521_assgn65217;
    reg [31:0] z2521_assgn2521;
    wire [31:0] a1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6525_assgn6525;
    reg [31:0] z6525_assgn65250;
    reg [31:0] z6525_assgn65251;
    reg [31:0] z6525_assgn65252;
    reg [31:0] z6525_assgn65253;
    reg [31:0] z6525_assgn65254;
    reg [31:0] z6525_assgn65255;
    reg [31:0] z6525_assgn65256;
    reg [31:0] z6525_assgn65257;
    reg [31:0] z2523_assgn2523;
    wire [31:0] a0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6529_assgn6529;
    reg [31:0] z6529_assgn65290;
    reg [31:0] z6529_assgn65291;
    reg [31:0] z6529_assgn65292;
    reg [31:0] z6529_assgn65293;
    reg [31:0] z6529_assgn65294;
    reg [31:0] z6529_assgn65295;
    reg [31:0] z6529_assgn65296;
    reg [31:0] z6529_assgn65297;
    reg [31:0] z2525_assgn2525;
    wire [31:0] a1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6533_assgn6533;
    reg [31:0] z6533_assgn65330;
    reg [31:0] z6533_assgn65331;
    reg [31:0] z6533_assgn65332;
    reg [31:0] z6533_assgn65333;
    reg [31:0] z6533_assgn65334;
    reg [31:0] z6533_assgn65335;
    reg [31:0] z6533_assgn65336;
    reg [31:0] z6533_assgn65337;
    reg [31:0] z2527_assgn2527;
    wire [31:0] b0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6537_assgn6537;
    reg [31:0] z6537_assgn65370;
    reg [31:0] z6537_assgn65371;
    reg [31:0] z6537_assgn65372;
    reg [31:0] z6537_assgn65373;
    reg [31:0] z6537_assgn65374;
    reg [31:0] z6537_assgn65375;
    reg [31:0] z6537_assgn65376;
    reg [31:0] z6537_assgn65377;
    reg [31:0] z2529_assgn2529;
    wire [31:0] b1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6541_assgn6541;
    reg [31:0] z6541_assgn65410;
    reg [31:0] z6541_assgn65411;
    reg [31:0] z6541_assgn65412;
    reg [31:0] z6541_assgn65413;
    reg [31:0] z6541_assgn65414;
    reg [31:0] z2531_assgn2531;
    wire [31:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6545_assgn6545;
    reg [31:0] z6545_assgn65450;
    reg [31:0] z6545_assgn65451;
    reg [31:0] z6545_assgn65452;
    reg [31:0] z6545_assgn65453;
    reg [31:0] z6545_assgn65454;
    reg [31:0] z2533_assgn2533;
    wire [31:0] c1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6549_assgn6549;
    reg [31:0] z6549_assgn65490;
    reg [31:0] z6549_assgn65491;
    reg [31:0] z6549_assgn65492;
    reg [31:0] z6549_assgn65493;
    reg [31:0] z6549_assgn65494;
    reg [31:0] z2535_assgn2535;
    wire [31:0] c0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6553_assgn6553;
    reg [31:0] z6553_assgn65530;
    reg [31:0] z6553_assgn65531;
    reg [31:0] z6553_assgn65532;
    reg [31:0] z6553_assgn65533;
    reg [31:0] z6553_assgn65534;
    reg [31:0] z2537_assgn2537;
    wire [31:0] c1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6557_assgn6557;
    reg [31:0] z6557_assgn65570;
    reg [31:0] z6557_assgn65571;
    reg [31:0] z6557_assgn65572;
    reg [31:0] z6557_assgn65573;
    reg [31:0] z6557_assgn65574;
    reg [31:0] z2539_assgn2539;
    wire [31:0] d0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6561_assgn6561;
    reg [31:0] z6561_assgn65610;
    reg [31:0] z6561_assgn65611;
    reg [31:0] z6561_assgn65612;
    reg [31:0] z6561_assgn65613;
    reg [31:0] z6561_assgn65614;
    reg [31:0] z2541_assgn2541;
    wire [31:0] d1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] c0_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] d0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] c1_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] d1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] cxord_1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6573_assgn6573;
    reg [31:0] z6573_assgn65730;
    reg [31:0] z6573_assgn65731;
    reg [31:0] z6573_assgn65732;
    reg [31:0] z6573_assgn65733;
    reg [31:0] z6573_assgn65734;
    reg [31:0] z6573_assgn65735;
    reg [31:0] z2551_assgn2551;
    wire [31:0] r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6581_assgn6581;
    reg [31:0] z6581_assgn65810;
    reg [31:0] z2557_assgn2557;
    wire [31:0] u0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6585_assgn6585;
    reg [31:0] z6585_assgn65850;
    reg [31:0] z2559_assgn2559;
    wire [31:0] u1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] cxord_0_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] r0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] cxord_1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] v1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6593_assgn6593;
    reg [31:0] z6593_assgn65930;
    reg [31:0] z2565_assgn2565;
    wire [31:0] p0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] e0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6603_assgn6603;
    reg [31:0] z6603_assgn66030;
    reg [31:0] z2573_assgn2573;
    wire [31:0] p2_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] e1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6613_assgn6613;
    reg [31:0] z6613_assgn66130;
    reg [31:0] z6613_assgn66131;
    reg [31:0] z6613_assgn66132;
    reg [31:0] z6613_assgn66133;
    reg [31:0] z6613_assgn66134;
    reg [31:0] z6613_assgn66135;
    reg [31:0] z2581_assgn2581;
    wire [31:0] r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6621_assgn6621;
    reg [31:0] z6621_assgn66210;
    reg [31:0] z2587_assgn2587;
    wire [31:0] u0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6625_assgn6625;
    reg [31:0] z6625_assgn66250;
    reg [31:0] z2589_assgn2589;
    wire [31:0] u1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6629_assgn6629;
    reg [31:0] z6629_assgn66290;
    reg [31:0] z2592_assgn2592;
    reg [31:0] r0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6633_assgn6633;
    reg [31:0] z6633_assgn66330;
    reg [31:0] z2594_assgn2594;
    wire [31:0] v1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6637_assgn6637;
    reg [31:0] z6637_assgn66370;
    reg [31:0] z6637_assgn66371;
    reg [31:0] z2595_assgn2595;
    wire [31:0] p0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6647_assgn6647;
    reg [31:0] z6647_assgn66470;
    reg [31:0] z6647_assgn66471;
    reg [31:0] z2603_assgn2603;
    wire [31:0] p2_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6661_assgn6661;
    reg [31:0] z6661_assgn66610;
    reg [31:0] z6661_assgn66611;
    reg [31:0] z6661_assgn66612;
    reg [31:0] z6661_assgn66613;
    reg [31:0] z6661_assgn66614;
    reg [31:0] z6661_assgn66615;
    reg [31:0] z2615_assgn2615;
    wire [31:0] r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a0_neg_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a1_neg_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6669_assgn6669;
    reg [31:0] z6669_assgn66690;
    reg [31:0] z2621_assgn2621;
    wire [31:0] u0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6673_assgn6673;
    reg [31:0] z6673_assgn66730;
    reg [31:0] z2623_assgn2623;
    wire [31:0] u1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6677_assgn6677;
    reg [31:0] z6677_assgn66770;
    reg [31:0] z2626_assgn2626;
    reg [31:0] r0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] v0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6681_assgn6681;
    reg [31:0] z6681_assgn66810;
    reg [31:0] z2628_assgn2628;
    wire [31:0] v1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6685_assgn6685;
    reg [31:0] z6685_assgn66850;
    reg [31:0] z6685_assgn66851;
    reg [31:0] z2629_assgn2629;
    wire [31:0] p0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] v1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] u0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] p1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p01_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6695_assgn6695;
    reg [31:0] z6695_assgn66950;
    reg [31:0] z6695_assgn66951;
    reg [31:0] z2637_assgn2637;
    wire [31:0] p2_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] v0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] u1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] p3_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p23_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p2_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] q1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6709_assgn6709;
    reg [31:0] z6709_assgn67090;
    reg [31:0] z6709_assgn67091;
    reg [31:0] z6709_assgn67092;
    reg [31:0] z6709_assgn67093;
    reg [31:0] z6709_assgn67094;
    reg [31:0] z6709_assgn67095;
    reg [31:0] z6709_assgn67096;
    reg [31:0] z6709_assgn67097;
    reg [31:0] z6709_assgn67098;
    reg [31:0] z2649_assgn2649;
    wire [31:0] p1ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z6713_assgn6713;
    reg [31:0] z6713_assgn67130;
    reg [31:0] z6713_assgn67131;
    reg [31:0] z6713_assgn67132;
    reg [31:0] z6713_assgn67133;
    reg [31:0] z6713_assgn67134;
    reg [31:0] z6713_assgn67135;
    reg [31:0] z6713_assgn67136;
    reg [31:0] z6713_assgn67137;
    reg [31:0] z6713_assgn67138;
    reg [31:0] z2651_assgn2651;
    wire [31:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q0_0_G16_mul2_G256_inv0;
    wire [31:0] q1_0_G16_mul2_G256_inv0;
    wire [31:0] q0_G16_mul2_G256_inv0;
    wire [31:0] q1_G16_mul2_G256_inv0;
    wire [31:0] z6725_assgn6725;
    reg [31:0] z6725_assgn67250;
    reg [31:0] z6725_assgn67251;
    reg [31:0] z6725_assgn67252;
    reg [31:0] z6725_assgn67253;
    reg [31:0] z6725_assgn67254;
    reg [31:0] z6725_assgn67255;
    reg [31:0] z6725_assgn67256;
    reg [31:0] z6725_assgn67257;
    reg [31:0] z6725_assgn67258;
    reg [31:0] z2661_assgn2661;
    wire [31:0] p0ls2_G16_mul2_G256_inv0;
    wire [31:0] z6729_assgn6729;
    reg [31:0] z6729_assgn67290;
    reg [31:0] z6729_assgn67291;
    reg [31:0] z6729_assgn67292;
    reg [31:0] z6729_assgn67293;
    reg [31:0] z6729_assgn67294;
    reg [31:0] z6729_assgn67295;
    reg [31:0] z6729_assgn67296;
    reg [31:0] z6729_assgn67297;
    reg [31:0] z6729_assgn67298;
    reg [31:0] z2663_assgn2663;
    wire [31:0] p1ls2_G16_mul2_G256_inv0;
    wire [31:0] q0_G256_inv0;
    wire [31:0] q1_G256_inv0;
    wire [31:0] z6737_assgn6737;
    reg [31:0] z6737_assgn67370;
    reg [31:0] z6737_assgn67371;
    reg [31:0] z6737_assgn67372;
    reg [31:0] z6737_assgn67373;
    reg [31:0] z6737_assgn67374;
    reg [31:0] z6737_assgn67375;
    reg [31:0] z6737_assgn67376;
    reg [31:0] z6737_assgn67377;
    reg [31:0] z2669_assgn2669;
    wire [31:0] p0ls4_G256_inv0;
    wire [31:0] z6741_assgn6741;
    reg [31:0] z6741_assgn67410;
    reg [31:0] z6741_assgn67411;
    reg [31:0] z6741_assgn67412;
    reg [31:0] z6741_assgn67413;
    reg [31:0] z6741_assgn67414;
    reg [31:0] z6741_assgn67415;
    reg [31:0] z6741_assgn67416;
    reg [31:0] z6741_assgn67417;
    reg [31:0] z2671_assgn2671;
    wire [31:0] p1ls4_G256_inv0;
    wire [31:0] t4;
    wire [31:0] t5;
    wire [31:0] z6749_assgn6749;
    reg [31:0] z6749_assgn67490;
    reg [31:0] z6749_assgn67491;
    reg [31:0] z6749_assgn67492;
    reg [31:0] z6749_assgn67493;
    reg [31:0] z6749_assgn67494;
    reg [31:0] z6749_assgn67495;
    reg [31:0] z6749_assgn67496;
    reg [31:0] z6749_assgn67497;
    reg [31:0] z6749_assgn67498;
    reg [31:0] y_G256_newbasis1;
    wire [31:0] tempy1_G256_newbasis1;
    wire [31:0] z6753_assgn6753;
    reg [31:0] z6753_assgn67530;
    reg [31:0] z6753_assgn67531;
    reg [31:0] z6753_assgn67532;
    reg [31:0] z6753_assgn67533;
    reg [31:0] z6753_assgn67534;
    reg [31:0] z6753_assgn67535;
    reg [31:0] z6753_assgn67536;
    reg [31:0] z6753_assgn67537;
    reg [31:0] z6753_assgn67538;
    reg [31:0] z2681_assgn2681;
    wire [31:0] cond1_G256_newbasis1;
    wire [31:0] negCond1_G256_newbasis1;
    wire [31:0] yxorb1_G256_newbasis1;
    wire [31:0] ny1_G256_newbasis1;
    wire [31:0] tempyIntoNegCond1_G256_newbasis1;
    wire [31:0] y1_G256_newbasis1;
    wire [31:0] z6767_assgn6767;
    reg [31:0] z6767_assgn67670;
    reg [31:0] z6767_assgn67671;
    reg [31:0] z6767_assgn67672;
    reg [31:0] z6767_assgn67673;
    reg [31:0] z6767_assgn67674;
    reg [31:0] z6767_assgn67675;
    reg [31:0] z6767_assgn67676;
    reg [31:0] z6767_assgn67677;
    reg [31:0] z6767_assgn67678;
    reg [31:0] z2693_assgn2693;
    wire [31:0] x1_G256_newbasis1;
    wire [31:0] tempy2_G256_newbasis1;
    wire [31:0] z6773_assgn6773;
    reg [31:0] z6773_assgn67730;
    reg [31:0] z6773_assgn67731;
    reg [31:0] z6773_assgn67732;
    reg [31:0] z6773_assgn67733;
    reg [31:0] z6773_assgn67734;
    reg [31:0] z6773_assgn67735;
    reg [31:0] z6773_assgn67736;
    reg [31:0] z6773_assgn67737;
    reg [31:0] z6773_assgn67738;
    reg [31:0] z2697_assgn2697;
    wire [31:0] cond2_G256_newbasis1;
    wire [31:0] negCond2_G256_newbasis1;
    wire [31:0] z6779_assgn6779;
    reg [31:0] z6779_assgn67790;
    reg [31:0] z6779_assgn67791;
    reg [31:0] z6779_assgn67792;
    reg [31:0] z6779_assgn67793;
    reg [31:0] z6779_assgn67794;
    reg [31:0] z6779_assgn67795;
    reg [31:0] z6779_assgn67796;
    reg [31:0] z6779_assgn67797;
    reg [31:0] z6779_assgn67798;
    reg [31:0] z2701_assgn2701;
    wire [31:0] yxorb2_G256_newbasis1;
    wire [31:0] ny2_G256_newbasis1;
    wire [31:0] tempyIntoNegCond2_G256_newbasis1;
    wire [31:0] y2_G256_newbasis1;
    wire [31:0] z6789_assgn6789;
    reg [31:0] z6789_assgn67890;
    reg [31:0] z6789_assgn67891;
    reg [31:0] z6789_assgn67892;
    reg [31:0] z6789_assgn67893;
    reg [31:0] z6789_assgn67894;
    reg [31:0] z6789_assgn67895;
    reg [31:0] z6789_assgn67896;
    reg [31:0] z6789_assgn67897;
    reg [31:0] z6789_assgn67898;
    reg [31:0] z2709_assgn2709;
    wire [31:0] x2_G256_newbasis1;
    wire [31:0] tempy3_G256_newbasis1;
    wire [31:0] z6795_assgn6795;
    reg [31:0] z6795_assgn67950;
    reg [31:0] z6795_assgn67951;
    reg [31:0] z6795_assgn67952;
    reg [31:0] z6795_assgn67953;
    reg [31:0] z6795_assgn67954;
    reg [31:0] z6795_assgn67955;
    reg [31:0] z6795_assgn67956;
    reg [31:0] z6795_assgn67957;
    reg [31:0] z6795_assgn67958;
    reg [31:0] z2713_assgn2713;
    wire [31:0] cond3_G256_newbasis1;
    wire [31:0] negCond3_G256_newbasis1;
    wire [31:0] z6801_assgn6801;
    reg [31:0] z6801_assgn68010;
    reg [31:0] z6801_assgn68011;
    reg [31:0] z6801_assgn68012;
    reg [31:0] z6801_assgn68013;
    reg [31:0] z6801_assgn68014;
    reg [31:0] z6801_assgn68015;
    reg [31:0] z6801_assgn68016;
    reg [31:0] z6801_assgn68017;
    reg [31:0] z2717_assgn2717;
    wire [31:0] yxorb3_G256_newbasis1;
    wire [31:0] ny3_G256_newbasis1;
    wire [31:0] tempyIntoNegCond3_G256_newbasis1;
    wire [31:0] y3_G256_newbasis1;
    wire [31:0] z6811_assgn6811;
    reg [31:0] z6811_assgn68110;
    reg [31:0] z6811_assgn68111;
    reg [31:0] z6811_assgn68112;
    reg [31:0] z6811_assgn68113;
    reg [31:0] z6811_assgn68114;
    reg [31:0] z6811_assgn68115;
    reg [31:0] z6811_assgn68116;
    reg [31:0] z6811_assgn68117;
    reg [31:0] z6811_assgn68118;
    reg [31:0] z2725_assgn2725;
    wire [31:0] x3_G256_newbasis1;
    wire [31:0] tempy4_G256_newbasis1;
    wire [31:0] z6817_assgn6817;
    reg [31:0] z6817_assgn68170;
    reg [31:0] z6817_assgn68171;
    reg [31:0] z6817_assgn68172;
    reg [31:0] z6817_assgn68173;
    reg [31:0] z6817_assgn68174;
    reg [31:0] z6817_assgn68175;
    reg [31:0] z6817_assgn68176;
    reg [31:0] z6817_assgn68177;
    reg [31:0] z6817_assgn68178;
    reg [31:0] z2729_assgn2729;
    wire [31:0] cond4_G256_newbasis1;
    wire [31:0] negCond4_G256_newbasis1;
    wire [31:0] yxorb4_G256_newbasis1;
    wire [31:0] ny4_G256_newbasis1;
    wire [31:0] tempyIntoNegCond4_G256_newbasis1;
    wire [31:0] y4_G256_newbasis1;
    wire [31:0] z6831_assgn6831;
    reg [31:0] z6831_assgn68310;
    reg [31:0] z6831_assgn68311;
    reg [31:0] z6831_assgn68312;
    reg [31:0] z6831_assgn68313;
    reg [31:0] z6831_assgn68314;
    reg [31:0] z6831_assgn68315;
    reg [31:0] z6831_assgn68316;
    reg [31:0] z6831_assgn68317;
    reg [31:0] z6831_assgn68318;
    reg [31:0] z2741_assgn2741;
    wire [31:0] x4_G256_newbasis1;
    wire [31:0] tempy5_G256_newbasis1;
    wire [31:0] z6837_assgn6837;
    reg [31:0] z6837_assgn68370;
    reg [31:0] z6837_assgn68371;
    reg [31:0] z6837_assgn68372;
    reg [31:0] z6837_assgn68373;
    reg [31:0] z6837_assgn68374;
    reg [31:0] z6837_assgn68375;
    reg [31:0] z6837_assgn68376;
    reg [31:0] z6837_assgn68377;
    reg [31:0] z6837_assgn68378;
    reg [31:0] z2745_assgn2745;
    wire [31:0] cond5_G256_newbasis1;
    wire [31:0] negCond5_G256_newbasis1;
    wire [31:0] yxorb5_G256_newbasis1;
    wire [31:0] ny5_G256_newbasis1;
    wire [31:0] tempyIntoNegCond5_G256_newbasis1;
    wire [31:0] y5_G256_newbasis1;
    wire [31:0] z6851_assgn6851;
    reg [31:0] z6851_assgn68510;
    reg [31:0] z6851_assgn68511;
    reg [31:0] z6851_assgn68512;
    reg [31:0] z6851_assgn68513;
    reg [31:0] z6851_assgn68514;
    reg [31:0] z6851_assgn68515;
    reg [31:0] z6851_assgn68516;
    reg [31:0] z6851_assgn68517;
    reg [31:0] z6851_assgn68518;
    reg [31:0] z2757_assgn2757;
    wire [31:0] x5_G256_newbasis1;
    wire [31:0] tempy6_G256_newbasis1;
    wire [31:0] z6857_assgn6857;
    reg [31:0] z6857_assgn68570;
    reg [31:0] z6857_assgn68571;
    reg [31:0] z6857_assgn68572;
    reg [31:0] z6857_assgn68573;
    reg [31:0] z6857_assgn68574;
    reg [31:0] z6857_assgn68575;
    reg [31:0] z6857_assgn68576;
    reg [31:0] z6857_assgn68577;
    reg [31:0] z6857_assgn68578;
    reg [31:0] z2761_assgn2761;
    wire [31:0] cond6_G256_newbasis1;
    wire [31:0] negCond6_G256_newbasis1;
    wire [31:0] yxorb6_G256_newbasis1;
    wire [31:0] ny6_G256_newbasis1;
    wire [31:0] tempyIntoNegCond6_G256_newbasis1;
    wire [31:0] y6_G256_newbasis1;
    wire [31:0] z6871_assgn6871;
    reg [31:0] z6871_assgn68710;
    reg [31:0] z6871_assgn68711;
    reg [31:0] z6871_assgn68712;
    reg [31:0] z6871_assgn68713;
    reg [31:0] z6871_assgn68714;
    reg [31:0] z6871_assgn68715;
    reg [31:0] z6871_assgn68716;
    reg [31:0] z6871_assgn68717;
    reg [31:0] z6871_assgn68718;
    reg [31:0] z2773_assgn2773;
    wire [31:0] x6_G256_newbasis1;
    wire [31:0] tempy7_G256_newbasis1;
    wire [31:0] z6877_assgn6877;
    reg [31:0] z6877_assgn68770;
    reg [31:0] z6877_assgn68771;
    reg [31:0] z6877_assgn68772;
    reg [31:0] z6877_assgn68773;
    reg [31:0] z6877_assgn68774;
    reg [31:0] z6877_assgn68775;
    reg [31:0] z6877_assgn68776;
    reg [31:0] z6877_assgn68777;
    reg [31:0] z6877_assgn68778;
    reg [31:0] z2777_assgn2777;
    wire [31:0] cond7_G256_newbasis1;
    wire [31:0] negCond7_G256_newbasis1;
    wire [31:0] yxorb7_G256_newbasis1;
    wire [31:0] ny7_G256_newbasis1;
    wire [31:0] tempyIntoNegCond7_G256_newbasis1;
    wire [31:0] y7_G256_newbasis1;
    wire [31:0] z6891_assgn6891;
    reg [31:0] z6891_assgn68910;
    reg [31:0] z6891_assgn68911;
    reg [31:0] z6891_assgn68912;
    reg [31:0] z6891_assgn68913;
    reg [31:0] z6891_assgn68914;
    reg [31:0] z6891_assgn68915;
    reg [31:0] z6891_assgn68916;
    reg [31:0] z6891_assgn68917;
    reg [31:0] z6891_assgn68918;
    reg [31:0] z2789_assgn2789;
    wire [31:0] x7_G256_newbasis1;
    wire [31:0] tempy8_G256_newbasis1;
    wire [31:0] z6897_assgn6897;
    reg [31:0] z6897_assgn68970;
    reg [31:0] z6897_assgn68971;
    reg [31:0] z6897_assgn68972;
    reg [31:0] z6897_assgn68973;
    reg [31:0] z6897_assgn68974;
    reg [31:0] z6897_assgn68975;
    reg [31:0] z6897_assgn68976;
    reg [31:0] z6897_assgn68977;
    reg [31:0] z6897_assgn68978;
    reg [31:0] z2793_assgn2793;
    wire [31:0] cond8_G256_newbasis1;
    wire [31:0] negCond8_G256_newbasis1;
    wire [31:0] yxorb8_G256_newbasis1;
    wire [31:0] ny8_G256_newbasis1;
    wire [31:0] tempyIntoNegCond8_G256_newbasis1;
    wire [31:0] y8_G256_newbasis1;
    wire [31:0] z6911_assgn6911;
    reg [31:0] z6911_assgn69110;
    reg [31:0] z6911_assgn69111;
    reg [31:0] z6911_assgn69112;
    reg [31:0] z6911_assgn69113;
    reg [31:0] z6911_assgn69114;
    reg [31:0] z6911_assgn69115;
    reg [31:0] z6911_assgn69116;
    reg [31:0] z6911_assgn69117;
    reg [31:0] z6911_assgn69118;
    reg [31:0] z2805_assgn2805;
    wire [31:0] x8_G256_newbasis1;
    wire [31:0] t6;
    wire [31:0] z6917_assgn6917;
    reg [31:0] z6917_assgn69170;
    reg [31:0] z6917_assgn69171;
    reg [31:0] z6917_assgn69172;
    reg [31:0] z6917_assgn69173;
    reg [31:0] z6917_assgn69174;
    reg [31:0] z6917_assgn69175;
    reg [31:0] z6917_assgn69176;
    reg [31:0] z6917_assgn69177;
    reg [31:0] z6917_assgn69178;
    reg [31:0] z_y_G256_newbasis1;
    wire [31:0] z_tempy1_G256_newbasis1;
    wire [31:0] z6921_assgn6921;
    reg [31:0] z6921_assgn69210;
    reg [31:0] z6921_assgn69211;
    reg [31:0] z6921_assgn69212;
    reg [31:0] z6921_assgn69213;
    reg [31:0] z6921_assgn69214;
    reg [31:0] z6921_assgn69215;
    reg [31:0] z6921_assgn69216;
    reg [31:0] z6921_assgn69217;
    reg [31:0] z6921_assgn69218;
    reg [31:0] z2813_assgn2813;
    wire [31:0] z_cond1_G256_newbasis1;
    wire [31:0] z_negCond1_G256_newbasis1;
    wire [31:0] z_yxorb1_G256_newbasis1;
    wire [31:0] z_ny1_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond1_G256_newbasis1;
    wire [31:0] z_y1_G256_newbasis1;
    wire [31:0] z6935_assgn6935;
    reg [31:0] z6935_assgn69350;
    reg [31:0] z6935_assgn69351;
    reg [31:0] z6935_assgn69352;
    reg [31:0] z6935_assgn69353;
    reg [31:0] z6935_assgn69354;
    reg [31:0] z6935_assgn69355;
    reg [31:0] z6935_assgn69356;
    reg [31:0] z6935_assgn69357;
    reg [31:0] z6935_assgn69358;
    reg [31:0] z2825_assgn2825;
    wire [31:0] z_x1_G256_newbasis1;
    wire [31:0] z_tempy2_G256_newbasis1;
    wire [31:0] z6941_assgn6941;
    reg [31:0] z6941_assgn69410;
    reg [31:0] z6941_assgn69411;
    reg [31:0] z6941_assgn69412;
    reg [31:0] z6941_assgn69413;
    reg [31:0] z6941_assgn69414;
    reg [31:0] z6941_assgn69415;
    reg [31:0] z6941_assgn69416;
    reg [31:0] z6941_assgn69417;
    reg [31:0] z6941_assgn69418;
    reg [31:0] z2829_assgn2829;
    wire [31:0] z_cond2_G256_newbasis1;
    wire [31:0] z_negCond2_G256_newbasis1;
    wire [31:0] z6947_assgn6947;
    reg [31:0] z6947_assgn69470;
    reg [31:0] z6947_assgn69471;
    reg [31:0] z6947_assgn69472;
    reg [31:0] z6947_assgn69473;
    reg [31:0] z6947_assgn69474;
    reg [31:0] z6947_assgn69475;
    reg [31:0] z6947_assgn69476;
    reg [31:0] z6947_assgn69477;
    reg [31:0] z6947_assgn69478;
    reg [31:0] z2833_assgn2833;
    wire [31:0] z_yxorb2_G256_newbasis1;
    wire [31:0] z_ny2_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond2_G256_newbasis1;
    wire [31:0] z_y2_G256_newbasis1;
    wire [31:0] z6957_assgn6957;
    reg [31:0] z6957_assgn69570;
    reg [31:0] z6957_assgn69571;
    reg [31:0] z6957_assgn69572;
    reg [31:0] z6957_assgn69573;
    reg [31:0] z6957_assgn69574;
    reg [31:0] z6957_assgn69575;
    reg [31:0] z6957_assgn69576;
    reg [31:0] z6957_assgn69577;
    reg [31:0] z6957_assgn69578;
    reg [31:0] z2841_assgn2841;
    wire [31:0] z_x2_G256_newbasis1;
    wire [31:0] z_tempy3_G256_newbasis1;
    wire [31:0] z6963_assgn6963;
    reg [31:0] z6963_assgn69630;
    reg [31:0] z6963_assgn69631;
    reg [31:0] z6963_assgn69632;
    reg [31:0] z6963_assgn69633;
    reg [31:0] z6963_assgn69634;
    reg [31:0] z6963_assgn69635;
    reg [31:0] z6963_assgn69636;
    reg [31:0] z6963_assgn69637;
    reg [31:0] z6963_assgn69638;
    reg [31:0] z2845_assgn2845;
    wire [31:0] z_cond3_G256_newbasis1;
    wire [31:0] z_negCond3_G256_newbasis1;
    wire [31:0] z6969_assgn6969;
    reg [31:0] z6969_assgn69690;
    reg [31:0] z6969_assgn69691;
    reg [31:0] z6969_assgn69692;
    reg [31:0] z6969_assgn69693;
    reg [31:0] z6969_assgn69694;
    reg [31:0] z6969_assgn69695;
    reg [31:0] z6969_assgn69696;
    reg [31:0] z6969_assgn69697;
    reg [31:0] z2849_assgn2849;
    wire [31:0] z_yxorb3_G256_newbasis1;
    wire [31:0] z_ny3_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond3_G256_newbasis1;
    wire [31:0] z_y3_G256_newbasis1;
    wire [31:0] z6979_assgn6979;
    reg [31:0] z6979_assgn69790;
    reg [31:0] z6979_assgn69791;
    reg [31:0] z6979_assgn69792;
    reg [31:0] z6979_assgn69793;
    reg [31:0] z6979_assgn69794;
    reg [31:0] z6979_assgn69795;
    reg [31:0] z6979_assgn69796;
    reg [31:0] z6979_assgn69797;
    reg [31:0] z6979_assgn69798;
    reg [31:0] z2857_assgn2857;
    wire [31:0] z_x3_G256_newbasis1;
    wire [31:0] z_tempy4_G256_newbasis1;
    wire [31:0] z6985_assgn6985;
    reg [31:0] z6985_assgn69850;
    reg [31:0] z6985_assgn69851;
    reg [31:0] z6985_assgn69852;
    reg [31:0] z6985_assgn69853;
    reg [31:0] z6985_assgn69854;
    reg [31:0] z6985_assgn69855;
    reg [31:0] z6985_assgn69856;
    reg [31:0] z6985_assgn69857;
    reg [31:0] z6985_assgn69858;
    reg [31:0] z2861_assgn2861;
    wire [31:0] z_cond4_G256_newbasis1;
    wire [31:0] z_negCond4_G256_newbasis1;
    wire [31:0] z_yxorb4_G256_newbasis1;
    wire [31:0] z_ny4_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond4_G256_newbasis1;
    wire [31:0] z_y4_G256_newbasis1;
    wire [31:0] z6999_assgn6999;
    reg [31:0] z6999_assgn69990;
    reg [31:0] z6999_assgn69991;
    reg [31:0] z6999_assgn69992;
    reg [31:0] z6999_assgn69993;
    reg [31:0] z6999_assgn69994;
    reg [31:0] z6999_assgn69995;
    reg [31:0] z6999_assgn69996;
    reg [31:0] z6999_assgn69997;
    reg [31:0] z6999_assgn69998;
    reg [31:0] z2873_assgn2873;
    wire [31:0] z_x4_G256_newbasis1;
    wire [31:0] z_tempy5_G256_newbasis1;
    wire [31:0] z7005_assgn7005;
    reg [31:0] z7005_assgn70050;
    reg [31:0] z7005_assgn70051;
    reg [31:0] z7005_assgn70052;
    reg [31:0] z7005_assgn70053;
    reg [31:0] z7005_assgn70054;
    reg [31:0] z7005_assgn70055;
    reg [31:0] z7005_assgn70056;
    reg [31:0] z7005_assgn70057;
    reg [31:0] z7005_assgn70058;
    reg [31:0] z2877_assgn2877;
    wire [31:0] z_cond5_G256_newbasis1;
    wire [31:0] z_negCond5_G256_newbasis1;
    wire [31:0] z_yxorb5_G256_newbasis1;
    wire [31:0] z_ny5_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond5_G256_newbasis1;
    wire [31:0] z_y5_G256_newbasis1;
    wire [31:0] z7019_assgn7019;
    reg [31:0] z7019_assgn70190;
    reg [31:0] z7019_assgn70191;
    reg [31:0] z7019_assgn70192;
    reg [31:0] z7019_assgn70193;
    reg [31:0] z7019_assgn70194;
    reg [31:0] z7019_assgn70195;
    reg [31:0] z7019_assgn70196;
    reg [31:0] z7019_assgn70197;
    reg [31:0] z7019_assgn70198;
    reg [31:0] z2889_assgn2889;
    wire [31:0] z_x5_G256_newbasis1;
    wire [31:0] z_tempy6_G256_newbasis1;
    wire [31:0] z7025_assgn7025;
    reg [31:0] z7025_assgn70250;
    reg [31:0] z7025_assgn70251;
    reg [31:0] z7025_assgn70252;
    reg [31:0] z7025_assgn70253;
    reg [31:0] z7025_assgn70254;
    reg [31:0] z7025_assgn70255;
    reg [31:0] z7025_assgn70256;
    reg [31:0] z7025_assgn70257;
    reg [31:0] z7025_assgn70258;
    reg [31:0] z2893_assgn2893;
    wire [31:0] z_cond6_G256_newbasis1;
    wire [31:0] z_negCond6_G256_newbasis1;
    wire [31:0] z_yxorb6_G256_newbasis1;
    wire [31:0] z_ny6_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond6_G256_newbasis1;
    wire [31:0] z_y6_G256_newbasis1;
    wire [31:0] z7039_assgn7039;
    reg [31:0] z7039_assgn70390;
    reg [31:0] z7039_assgn70391;
    reg [31:0] z7039_assgn70392;
    reg [31:0] z7039_assgn70393;
    reg [31:0] z7039_assgn70394;
    reg [31:0] z7039_assgn70395;
    reg [31:0] z7039_assgn70396;
    reg [31:0] z7039_assgn70397;
    reg [31:0] z7039_assgn70398;
    reg [31:0] z2905_assgn2905;
    wire [31:0] z_x6_G256_newbasis1;
    wire [31:0] z_tempy7_G256_newbasis1;
    wire [31:0] z7045_assgn7045;
    reg [31:0] z7045_assgn70450;
    reg [31:0] z7045_assgn70451;
    reg [31:0] z7045_assgn70452;
    reg [31:0] z7045_assgn70453;
    reg [31:0] z7045_assgn70454;
    reg [31:0] z7045_assgn70455;
    reg [31:0] z7045_assgn70456;
    reg [31:0] z7045_assgn70457;
    reg [31:0] z7045_assgn70458;
    reg [31:0] z2909_assgn2909;
    wire [31:0] z_cond7_G256_newbasis1;
    wire [31:0] z_negCond7_G256_newbasis1;
    wire [31:0] z_yxorb7_G256_newbasis1;
    wire [31:0] z_ny7_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond7_G256_newbasis1;
    wire [31:0] z_y7_G256_newbasis1;
    wire [31:0] z7059_assgn7059;
    reg [31:0] z7059_assgn70590;
    reg [31:0] z7059_assgn70591;
    reg [31:0] z7059_assgn70592;
    reg [31:0] z7059_assgn70593;
    reg [31:0] z7059_assgn70594;
    reg [31:0] z7059_assgn70595;
    reg [31:0] z7059_assgn70596;
    reg [31:0] z7059_assgn70597;
    reg [31:0] z7059_assgn70598;
    reg [31:0] z2921_assgn2921;
    wire [31:0] z_x7_G256_newbasis1;
    wire [31:0] z_tempy8_G256_newbasis1;
    wire [31:0] z7065_assgn7065;
    reg [31:0] z7065_assgn70650;
    reg [31:0] z7065_assgn70651;
    reg [31:0] z7065_assgn70652;
    reg [31:0] z7065_assgn70653;
    reg [31:0] z7065_assgn70654;
    reg [31:0] z7065_assgn70655;
    reg [31:0] z7065_assgn70656;
    reg [31:0] z7065_assgn70657;
    reg [31:0] z7065_assgn70658;
    reg [31:0] z2925_assgn2925;
    wire [31:0] z_cond8_G256_newbasis1;
    wire [31:0] z_negCond8_G256_newbasis1;
    wire [31:0] z_yxorb8_G256_newbasis1;
    wire [31:0] z_ny8_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond8_G256_newbasis1;
    wire [31:0] z_y8_G256_newbasis1;
    wire [31:0] z7079_assgn7079;
    reg [31:0] z7079_assgn70790;
    reg [31:0] z7079_assgn70791;
    reg [31:0] z7079_assgn70792;
    reg [31:0] z7079_assgn70793;
    reg [31:0] z7079_assgn70794;
    reg [31:0] z7079_assgn70795;
    reg [31:0] z7079_assgn70796;
    reg [31:0] z7079_assgn70797;
    reg [31:0] z7079_assgn70798;
    reg [31:0] z2937_assgn2937;
    wire [31:0] z_x8_G256_newbasis1;
    wire [31:0] t7;

    assign z2945_assgn2945 = dec_99;
    assign z2947_assgn2947 = dec_88;
    assign z2949_assgn2949 = dec_45;
    assign z2951_assgn2951 = dec_158;
    assign z2953_assgn2953 = dec_11;
    assign z2955_assgn2955 = dec_220;
    assign z2957_assgn2957 = dec_36;
    assign dec_16_inp = dec_16;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign z2975_assgn2975 = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t0_inp = t0;
    assign t1_inp = t1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign r3_inp = r3;
    assign r4_inp = r4;
    assign r5_inp = r5;
    assign r6_inp = r6;
    assign r7_inp = r7;
    assign r8_inp = r8;
    assign z3037_assgn3037 = r9;
    assign z3039_assgn3039 = r10;
    assign z3041_assgn3041 = r11;
    assign z3043_assgn3043 = r12;
    assign z3045_assgn3045 = r13;
    assign z3047_assgn3047 = r14;
    assign z3049_assgn3049 = r15;
    assign z3051_assgn3051 = r16;
    assign z3053_assgn3053 = r17;
    assign z3055_assgn3055 = r18;
    assign z3057_assgn3057 = r19;
    assign z3059_assgn3059 = r20;
    assign z3061_assgn3061 = r21;
    assign z3063_assgn3063 = r22;
    assign z3065_assgn3065 = r23;
    assign z3067_assgn3067 = r24;
    assign z3069_assgn3069 = r25;
    assign z3071_assgn3071 = r26;
    assign z3073_assgn3073 = r27;
    assign z3075_assgn3075 = r28;
    assign z3077_assgn3077 = r29;
    assign z3079_assgn3079 = r30;
    assign z3081_assgn3081 = r31;
    assign z3083_assgn3083 = r32;
    assign z3085_assgn3085 = r33;
    assign z3087_assgn3087 = r34;
    assign z3089_assgn3089 = r35;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t0_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempyIntoNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempyIntoNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t0_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempyIntoNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempyIntoNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempyIntoNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempyIntoNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempyIntoNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempyIntoNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempyIntoNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempyIntoNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempyIntoNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempyIntoNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempyIntoNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempyIntoNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempyIntoNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0);
    assign z3219_assgn3219 = dec_1_inp;
    assign z3221_assgn3221 = x7_G256_newbasis0;
    assign x8_G256_newbasis0 = (z298_assgn298 >> z297_assgn297);
    assign t2 = y8_G256_newbasis0;
    assign z_y_G256_newbasis0 = dec_0_inp;
    assign z_tempy1_G256_newbasis0 = z_y_G256_newbasis0;
    assign z_cond1_G256_newbasis0 = (t1_inp & dec_1_inp);
    assign z_negCond1_G256_newbasis0 = !z_cond1_G256_newbasis0;
    assign z_yxorb1_G256_newbasis0 = (z_y_G256_newbasis0 ^ dec_255_inp);
    assign z_ny1_G256_newbasis0 = (z_cond1_G256_newbasis0 * z_yxorb1_G256_newbasis0);
    assign z_tempyIntoNegCond1_G256_newbasis0 = (z_tempy1_G256_newbasis0 * z_negCond1_G256_newbasis0);
    assign z_y1_G256_newbasis0 = (z_ny1_G256_newbasis0 + z_tempyIntoNegCond1_G256_newbasis0);
    assign z_x1_G256_newbasis0 = (t1_inp >> dec_1_inp);
    assign z_tempy2_G256_newbasis0 = z_y1_G256_newbasis0;
    assign z_cond2_G256_newbasis0 = (z_x1_G256_newbasis0 & dec_1_inp);
    assign z_negCond2_G256_newbasis0 = !z_cond2_G256_newbasis0;
    assign z_yxorb2_G256_newbasis0 = (z_y1_G256_newbasis0 ^ dec_169_inp);
    assign z_ny2_G256_newbasis0 = (z_cond2_G256_newbasis0 * z_yxorb2_G256_newbasis0);
    assign z_tempyIntoNegCond2_G256_newbasis0 = (z_tempy2_G256_newbasis0 * z_negCond2_G256_newbasis0);
    assign z_y2_G256_newbasis0 = (z_ny2_G256_newbasis0 + z_tempyIntoNegCond2_G256_newbasis0);
    assign z_x2_G256_newbasis0 = (z_x1_G256_newbasis0 >> dec_1_inp);
    assign z_tempy3_G256_newbasis0 = z_y2_G256_newbasis0;
    assign z_cond3_G256_newbasis0 = (z_x2_G256_newbasis0 & dec_1_inp);
    assign z_negCond3_G256_newbasis0 = !z_cond3_G256_newbasis0;
    assign z_yxorb3_G256_newbasis0 = (z_y2_G256_newbasis0 ^ dec_129_inp);
    assign z_ny3_G256_newbasis0 = (z_cond3_G256_newbasis0 * z_yxorb3_G256_newbasis0);
    assign z_tempyIntoNegCond3_G256_newbasis0 = (z_tempy3_G256_newbasis0 * z_negCond3_G256_newbasis0);
    assign z_y3_G256_newbasis0 = (z_ny3_G256_newbasis0 + z_tempyIntoNegCond3_G256_newbasis0);
    assign z_x3_G256_newbasis0 = (z_x2_G256_newbasis0 >> dec_1_inp);
    assign z_tempy4_G256_newbasis0 = z_y3_G256_newbasis0;
    assign z_cond4_G256_newbasis0 = (z_x3_G256_newbasis0 & dec_1_inp);
    assign z_negCond4_G256_newbasis0 = !z_cond4_G256_newbasis0;
    assign z_yxorb4_G256_newbasis0 = (z_y3_G256_newbasis0 ^ dec_9_inp);
    assign z_ny4_G256_newbasis0 = (z_cond4_G256_newbasis0 * z_yxorb4_G256_newbasis0);
    assign z_tempyIntoNegCond4_G256_newbasis0 = (z_tempy4_G256_newbasis0 * z_negCond4_G256_newbasis0);
    assign z_y4_G256_newbasis0 = (z_ny4_G256_newbasis0 + z_tempyIntoNegCond4_G256_newbasis0);
    assign z_x4_G256_newbasis0 = (z_x3_G256_newbasis0 >> dec_1_inp);
    assign z_tempy5_G256_newbasis0 = z_y4_G256_newbasis0;
    assign z_cond5_G256_newbasis0 = (z_x4_G256_newbasis0 & dec_1_inp);
    assign z_negCond5_G256_newbasis0 = !z_cond5_G256_newbasis0;
    assign z_yxorb5_G256_newbasis0 = (z_y4_G256_newbasis0 ^ dec_72_inp);
    assign z_ny5_G256_newbasis0 = (z_cond5_G256_newbasis0 * z_yxorb5_G256_newbasis0);
    assign z_tempyIntoNegCond5_G256_newbasis0 = (z_tempy5_G256_newbasis0 * z_negCond5_G256_newbasis0);
    assign z_y5_G256_newbasis0 = (z_ny5_G256_newbasis0 + z_tempyIntoNegCond5_G256_newbasis0);
    assign z_x5_G256_newbasis0 = (z_x4_G256_newbasis0 >> dec_1_inp);
    assign z_tempy6_G256_newbasis0 = z_y5_G256_newbasis0;
    assign z_cond6_G256_newbasis0 = (z_x5_G256_newbasis0 & dec_1_inp);
    assign z_negCond6_G256_newbasis0 = !z_cond6_G256_newbasis0;
    assign z_yxorb6_G256_newbasis0 = (z_y5_G256_newbasis0 ^ dec_242_inp);
    assign z_ny6_G256_newbasis0 = (z_cond6_G256_newbasis0 * z_yxorb6_G256_newbasis0);
    assign z_tempyIntoNegCond6_G256_newbasis0 = (z_tempy6_G256_newbasis0 * z_negCond6_G256_newbasis0);
    assign z_y6_G256_newbasis0 = (z_ny6_G256_newbasis0 + z_tempyIntoNegCond6_G256_newbasis0);
    assign z_x6_G256_newbasis0 = (z_x5_G256_newbasis0 >> dec_1_inp);
    assign z_tempy7_G256_newbasis0 = z_y6_G256_newbasis0;
    assign z_cond7_G256_newbasis0 = (z_x6_G256_newbasis0 & dec_1_inp);
    assign z_negCond7_G256_newbasis0 = !z_cond7_G256_newbasis0;
    assign z_yxorb7_G256_newbasis0 = (z_y6_G256_newbasis0 ^ dec_243_inp);
    assign z_ny7_G256_newbasis0 = (z_cond7_G256_newbasis0 * z_yxorb7_G256_newbasis0);
    assign z_tempyIntoNegCond7_G256_newbasis0 = (z_tempy7_G256_newbasis0 * z_negCond7_G256_newbasis0);
    assign z_y7_G256_newbasis0 = (z_ny7_G256_newbasis0 + z_tempyIntoNegCond7_G256_newbasis0);
    assign z_x7_G256_newbasis0 = (z_x6_G256_newbasis0 >> dec_1_inp);
    assign z_tempy8_G256_newbasis0 = z_y7_G256_newbasis0;
    assign z_cond8_G256_newbasis0 = (z_x7_G256_newbasis0 & dec_1_inp);
    assign z_negCond8_G256_newbasis0 = !z_cond8_G256_newbasis0;
    assign z_yxorb8_G256_newbasis0 = (z_y7_G256_newbasis0 ^ dec_152_inp);
    assign z_ny8_G256_newbasis0 = (z_cond8_G256_newbasis0 * z_yxorb8_G256_newbasis0);
    assign z_tempyIntoNegCond8_G256_newbasis0 = (z_tempy8_G256_newbasis0 * z_negCond8_G256_newbasis0);
    assign z_y8_G256_newbasis0 = (z_ny8_G256_newbasis0 + z_tempyIntoNegCond8_G256_newbasis0);
    assign z3355_assgn3355 = dec_1_inp;
    assign z3357_assgn3357 = z_x7_G256_newbasis0;
    assign z_x8_G256_newbasis0 = (z430_assgn430 >> z429_assgn429);
    assign t3 = z_y8_G256_newbasis0;
    assign z3363_assgn3363 = t2;
    assign a0_0_G256_inv0 = (z434_assgn434 & dec_240_inp);
    assign z3367_assgn3367 = t3;
    assign a1_0_G256_inv0 = (z436_assgn436 & dec_240_inp);
    assign z3371_assgn3371 = z3_assgn3;
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> z437_assgn437);
    assign z3375_assgn3375 = z3_assgn3;
    assign a1_G256_inv0 = (a1_0_G256_inv0 >> z439_assgn439);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign b1_G256_inv0 = (t3 & dec_15_inp);
    assign z3383_assgn3383 = b0_G256_inv0;
    assign a0xorb0_G256_inv0 = (a0_G256_inv0_reg ^ z445_assgn445);
    assign z3387_assgn3387 = b1_G256_inv0;
    assign a1xorb1_G256_inv0 = (a1_G256_inv0_reg ^ z447_assgn447);
    assign z3391_assgn3391 = dec_12_inp;
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & z449_assgn449);
    assign z3395_assgn3395 = dec_12_inp;
    assign a1_0_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & z451_assgn451);
    assign z3399_assgn3399 = dec_2_inp;
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> z453_assgn453);
    assign z3403_assgn3403 = dec_2_inp;
    assign a1_G16_sq_scl0_G256_inv0 = (a1_0_G16_sq_scl0_G256_inv0 >> z455_assgn455);
    assign z3407_assgn3407 = dec_3_inp;
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & z457_assgn457);
    assign z3411_assgn3411 = dec_3_inp;
    assign b1_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & z459_assgn459);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign p1_0_G16_sq_scl0_G256_inv0 = (a1_G16_sq_scl0_G256_inv0 ^ b1_G16_sq_scl0_G256_inv0);
    assign z3419_assgn3419 = dec_2_inp;
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & z465_assgn465);
    assign z3423_assgn3423 = dec_2_inp;
    assign a1_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & z467_assgn467);
    assign z3427_assgn3427 = dec_1_inp;
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> z469_assgn469);
    assign z3431_assgn3431 = dec_1_inp;
    assign a1_G4_sq0_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq0_G16_sq_scl0_G256_inv0 >> z471_assgn471);
    assign z3435_assgn3435 = dec_1_inp;
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & z473_assgn473);
    assign z3439_assgn3439 = dec_1_inp;
    assign b1_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & z475_assgn475);
    assign z3443_assgn3443 = dec_1_inp;
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << z477_assgn477);
    assign z3447_assgn3447 = dec_1_inp;
    assign b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b1_G4_sq0_G16_sq_scl0_G256_inv0 << z479_assgn479);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign p1_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a1_G4_sq0_G16_sq_scl0_G256_inv0);
    assign z3455_assgn3455 = dec_2_inp;
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & z485_assgn485);
    assign z3459_assgn3459 = dec_2_inp;
    assign a1_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & z487_assgn487);
    assign z3463_assgn3463 = dec_1_inp;
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> z489_assgn489);
    assign z3467_assgn3467 = dec_1_inp;
    assign a1_G4_sq1_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq1_G16_sq_scl0_G256_inv0 >> z491_assgn491);
    assign z3471_assgn3471 = dec_1_inp;
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & z493_assgn493);
    assign z3475_assgn3475 = dec_1_inp;
    assign b1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & z495_assgn495);
    assign z3479_assgn3479 = dec_1_inp;
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << z497_assgn497);
    assign z3483_assgn3483 = dec_1_inp;
    assign b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G4_sq1_G16_sq_scl0_G256_inv0 << z499_assgn499);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign q1_0_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a1_G4_sq1_G16_sq_scl0_G256_inv0);
    assign z3491_assgn3491 = dec_2_inp;
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & z505_assgn505);
    assign z3495_assgn3495 = dec_2_inp;
    assign a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & z507_assgn507);
    assign z3499_assgn3499 = dec_1_inp;
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> z509_assgn509);
    assign z3503_assgn3503 = dec_1_inp;
    assign a1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> z511_assgn511);
    assign z3507_assgn3507 = dec_1_inp;
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & z513_assgn513);
    assign z3511_assgn3511 = dec_1_inp;
    assign b1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & z515_assgn515);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign q1_G4_scl_N20_G16_sq_scl0_G256_inv0 = a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign z3523_assgn3523 = dec_1_inp;
    assign p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p1_G4_scl_N20_G16_sq_scl0_G256_inv0 << z525_assgn525);
    assign z3527_assgn3527 = dec_1_inp;
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << z527_assgn527);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q1_G16_sq_scl0_G256_inv0 = (p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign z3535_assgn3535 = dec_2_inp;
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << z533_assgn533);
    assign z3539_assgn3539 = dec_2_inp;
    assign p1ls2_G16_sq_scl0_G256_inv0 = (p1_G16_sq_scl0_G256_inv0 << z535_assgn535);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign c1_G256_inv0 = (p1ls2_G16_sq_scl0_G256_inv0 | q1_G16_sq_scl0_G256_inv0);
    assign r00_G16_mul0_G256_inv0 = (z5_assgn5 % z1_assgn1);
    assign r10_G16_mul0_G256_inv0 = (z7_assgn7 % z1_assgn1);
    assign r20_G16_mul0_G256_inv0 = (z9_assgn9 % z1_assgn1);
    assign r30_G16_mul0_G256_inv0 = (z11_assgn11 % z1_assgn1);
    assign r40_G16_mul0_G256_inv0 = (z13_assgn13 % z1_assgn1);
    assign r50_G16_mul0_G256_inv0 = (z15_assgn15 % z1_assgn1);
    assign r60_G16_mul0_G256_inv0 = (z17_assgn17 % z1_assgn1);
    assign r70_G16_mul0_G256_inv0 = (z19_assgn19 % z1_assgn1);
    assign r80_G16_mul0_G256_inv0 = (z21_assgn21 % z1_assgn1);
    assign z3565_assgn3565 = dec_12_inp;
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & z559_assgn559);
    assign z3569_assgn3569 = dec_12_inp;
    assign a1_0_G16_mul0_G256_inv0 = (a1_G256_inv0 & z561_assgn561);
    assign z3573_assgn3573 = dec_2_inp;
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> z563_assgn563);
    assign z3577_assgn3577 = dec_2_inp;
    assign a1_G16_mul0_G256_inv0 = (a1_0_G16_mul0_G256_inv0 >> z565_assgn565);
    assign z3581_assgn3581 = dec_3_inp;
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & z567_assgn567);
    assign z3585_assgn3585 = dec_3_inp;
    assign b1_G16_mul0_G256_inv0 = (a1_G256_inv0 & z569_assgn569);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul0_G256_inv0 = (c1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign axorb_1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 ^ b1_G16_mul0_G256_inv0);
    assign cxord_1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 ^ d1_G16_mul0_G256_inv0);
    assign r00_G4_mul0_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % z3_assgn3);
    assign r10_G4_mul0_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % z3_assgn3);
    assign r20_G4_mul0_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % z3_assgn3);
    assign z3615_assgn3615 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & z597_assgn597);
    assign z3619_assgn3619 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & z599_assgn599);
    assign z3623_assgn3623 = dec_1_inp;
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> z601_assgn601);
    assign z3627_assgn3627 = dec_1_inp;
    assign a1_G4_mul0_G16_mul0_G256_inv0 = (a1_0_G4_mul0_G16_mul0_G256_inv0 >> z603_assgn603);
    assign z3631_assgn3631 = dec_1_inp;
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & z605_assgn605);
    assign z3635_assgn3635 = dec_1_inp;
    assign b1_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & z607_assgn607);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul0_G256_inv0 = (c1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0_reg ^ d0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign axorb_1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ b1_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0_reg ^ d1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign r0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0 = !axorb_0_G4_mul0_G16_mul0_G256_inv0;
    assign a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0 = !axorb_1_G4_mul0_G16_mul0_G256_inv0;
    assign z3665_assgn3665 = r0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    assign u0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0 & z635_assgn635);
    assign z3669_assgn3669 = r0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    assign u1_hpc20_G4_mul0_G16_mul0_G256_inv0 = (a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0 & z637_assgn637);
    assign v0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G4_mul0_G16_mul0_G256_inv0_reg ^ r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign v1_hpc20_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G4_mul0_G16_mul0_G256_inv0_reg ^ r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign z3677_assgn3677 = cxord_0_G4_mul0_G16_mul0_G256_inv0;
    assign p0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 & z643_assgn643);
    assign p1_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 & v1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p01_hpc20_G4_mul0_G16_mul0_G256_inv0 = (u0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul0_G256_inv0 = (p0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p01_hpc20_G4_mul0_G16_mul0_G256_inv0);
    assign z3687_assgn3687 = cxord_1_G4_mul0_G16_mul0_G256_inv0;
    assign p2_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0 & z651_assgn651);
    assign p3_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0 & v0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p23_hpc20_G4_mul0_G16_mul0_G256_inv0 = (u1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p3_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p23_hpc20_G4_mul0_G16_mul0_G256_inv0);
    assign r0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0 = !a0_G4_mul0_G16_mul0_G256_inv0;
    assign a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0 = !a1_G4_mul0_G16_mul0_G256_inv0;
    assign z3703_assgn3703 = r0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    assign u0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0 & z665_assgn665);
    assign z3707_assgn3707 = r0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    assign u1_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0 & z667_assgn667);
    assign z3711_assgn3711 = c0_G4_mul0_G16_mul0_G256_inv0;
    assign v0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (z670_assgn670 ^ r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign z3715_assgn3715 = c1_G4_mul0_G16_mul0_G256_inv0;
    assign v1_hpc21_G4_mul0_G16_mul0_G256_inv0 = (z672_assgn672 ^ r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign z3719_assgn3719 = c0_G4_mul0_G16_mul0_G256_inv0;
    assign p0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 & z673_assgn673);
    assign p1_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 & v1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p01_hpc21_G4_mul0_G16_mul0_G256_inv0 = (u0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (p0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p01_hpc21_G4_mul0_G16_mul0_G256_inv0);
    assign z3729_assgn3729 = c1_G4_mul0_G16_mul0_G256_inv0;
    assign p2_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 & z681_assgn681);
    assign p3_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 & v0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p23_hpc21_G4_mul0_G16_mul0_G256_inv0 = (u1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p3_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p23_hpc21_G4_mul0_G16_mul0_G256_inv0);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_G4_mul0_G16_mul0_G256_inv0 = (p1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign r0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0 = !b0_G4_mul0_G16_mul0_G256_inv0;
    assign a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0 = !b1_G4_mul0_G16_mul0_G256_inv0;
    assign z3749_assgn3749 = r0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    assign u0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0 & z699_assgn699);
    assign z3753_assgn3753 = r0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    assign u1_hpc22_G4_mul0_G16_mul0_G256_inv0 = (a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0 & z701_assgn701);
    assign z3757_assgn3757 = d0_G4_mul0_G16_mul0_G256_inv0;
    assign v0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (z704_assgn704 ^ r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign z3761_assgn3761 = d1_G4_mul0_G16_mul0_G256_inv0;
    assign v1_hpc22_G4_mul0_G16_mul0_G256_inv0 = (z706_assgn706 ^ r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign z3765_assgn3765 = d0_G4_mul0_G16_mul0_G256_inv0;
    assign p0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 & z707_assgn707);
    assign p1_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 & v1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p01_hpc22_G4_mul0_G16_mul0_G256_inv0 = (u0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (p0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p01_hpc22_G4_mul0_G16_mul0_G256_inv0);
    assign z3775_assgn3775 = d1_G4_mul0_G16_mul0_G256_inv0;
    assign p2_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0 & z715_assgn715);
    assign p3_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0 & v0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p23_hpc22_G4_mul0_G16_mul0_G256_inv0 = (u1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p3_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p23_hpc22_G4_mul0_G16_mul0_G256_inv0);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q1_G4_mul0_G16_mul0_G256_inv0 = (q1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign z3789_assgn3789 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul0_G256_inv0 = (p1_G4_mul0_G16_mul0_G256_inv0 << z727_assgn727);
    assign z3793_assgn3793 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << z729_assgn729);
    assign e0_G16_mul0_G256_inv0 = (p1ls1_G4_mul0_G16_mul0_G256_inv0 | q1_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign z3801_assgn3801 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & z735_assgn735);
    assign z3805_assgn3805 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z737_assgn737);
    assign z3809_assgn3809 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> z739_assgn739);
    assign z3813_assgn3813 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_0_G4_scl_N0_G16_mul0_G256_inv0 >> z741_assgn741);
    assign z3817_assgn3817 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & z743_assgn743);
    assign z3821_assgn3821 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z745_assgn745);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign p1_G4_scl_N0_G16_mul0_G256_inv0 = b1_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign q1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_G4_scl_N0_G16_mul0_G256_inv0 ^ b1_G4_scl_N0_G16_mul0_G256_inv0);
    assign z3833_assgn3833 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p1_G4_scl_N0_G16_mul0_G256_inv0 << z755_assgn755);
    assign z3837_assgn3837 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << z757_assgn757);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign e11_G16_mul0_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul0_G256_inv0 | q1_G4_scl_N0_G16_mul0_G256_inv0);
    assign r00_G4_mul1_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % z3_assgn3);
    assign r10_G4_mul1_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % z3_assgn3);
    assign r20_G4_mul1_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % z3_assgn3);
    assign z3851_assgn3851 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & z769_assgn769);
    assign z3855_assgn3855 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & z771_assgn771);
    assign z3859_assgn3859 = dec_1_inp;
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> z773_assgn773);
    assign z3863_assgn3863 = dec_1_inp;
    assign a1_G4_mul1_G16_mul0_G256_inv0 = (a1_0_G4_mul1_G16_mul0_G256_inv0 >> z775_assgn775);
    assign z3867_assgn3867 = dec_1_inp;
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & z777_assgn777);
    assign z3871_assgn3871 = dec_1_inp;
    assign b1_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & z779_assgn779);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul0_G256_inv0 = (c1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0_reg ^ d0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign axorb_1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ b1_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0_reg ^ d1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign r0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0 = !axorb_0_G4_mul1_G16_mul0_G256_inv0;
    assign a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0 = !axorb_1_G4_mul1_G16_mul0_G256_inv0;
    assign z3901_assgn3901 = r0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    assign u0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0 & z807_assgn807);
    assign z3905_assgn3905 = r0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    assign u1_hpc20_G4_mul1_G16_mul0_G256_inv0 = (a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0 & z809_assgn809);
    assign v0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (cxord_0_G4_mul1_G16_mul0_G256_inv0_reg ^ r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign v1_hpc20_G4_mul1_G16_mul0_G256_inv0 = (cxord_1_G4_mul1_G16_mul0_G256_inv0_reg ^ r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign z3913_assgn3913 = cxord_0_G4_mul1_G16_mul0_G256_inv0;
    assign p0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 & z815_assgn815);
    assign p1_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 & v1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p01_hpc20_G4_mul1_G16_mul0_G256_inv0 = (u0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul0_G256_inv0 = (p0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p01_hpc20_G4_mul1_G16_mul0_G256_inv0);
    assign z3923_assgn3923 = cxord_1_G4_mul1_G16_mul0_G256_inv0;
    assign p2_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0 & z823_assgn823);
    assign p3_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0 & v0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p23_hpc20_G4_mul1_G16_mul0_G256_inv0 = (u1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p3_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p23_hpc20_G4_mul1_G16_mul0_G256_inv0);
    assign r0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0 = !a0_G4_mul1_G16_mul0_G256_inv0;
    assign a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0 = !a1_G4_mul1_G16_mul0_G256_inv0;
    assign z3939_assgn3939 = r0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    assign u0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0 & z837_assgn837);
    assign z3943_assgn3943 = r0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    assign u1_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0 & z839_assgn839);
    assign z3947_assgn3947 = c0_G4_mul1_G16_mul0_G256_inv0;
    assign v0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (z842_assgn842 ^ r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign z3951_assgn3951 = c1_G4_mul1_G16_mul0_G256_inv0;
    assign v1_hpc21_G4_mul1_G16_mul0_G256_inv0 = (z844_assgn844 ^ r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign z3955_assgn3955 = c0_G4_mul1_G16_mul0_G256_inv0;
    assign p0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 & z845_assgn845);
    assign p1_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 & v1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p01_hpc21_G4_mul1_G16_mul0_G256_inv0 = (u0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (p0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p01_hpc21_G4_mul1_G16_mul0_G256_inv0);
    assign z3965_assgn3965 = c1_G4_mul1_G16_mul0_G256_inv0;
    assign p2_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 & z853_assgn853);
    assign p3_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 & v0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p23_hpc21_G4_mul1_G16_mul0_G256_inv0 = (u1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p3_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p23_hpc21_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_G4_mul1_G16_mul0_G256_inv0 = (p1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign r0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0 = !b0_G4_mul1_G16_mul0_G256_inv0;
    assign a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0 = !b1_G4_mul1_G16_mul0_G256_inv0;
    assign z3985_assgn3985 = r0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    assign u0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0 & z871_assgn871);
    assign z3989_assgn3989 = r0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    assign u1_hpc22_G4_mul1_G16_mul0_G256_inv0 = (a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0 & z873_assgn873);
    assign z3993_assgn3993 = d0_G4_mul1_G16_mul0_G256_inv0;
    assign v0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (z876_assgn876 ^ r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign z3997_assgn3997 = d1_G4_mul1_G16_mul0_G256_inv0;
    assign v1_hpc22_G4_mul1_G16_mul0_G256_inv0 = (z878_assgn878 ^ r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign z4001_assgn4001 = d0_G4_mul1_G16_mul0_G256_inv0;
    assign p0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 & z879_assgn879);
    assign p1_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 & v1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p01_hpc22_G4_mul1_G16_mul0_G256_inv0 = (u0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (p0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p01_hpc22_G4_mul1_G16_mul0_G256_inv0);
    assign z4011_assgn4011 = d1_G4_mul1_G16_mul0_G256_inv0;
    assign p2_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0 & z887_assgn887);
    assign p3_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0 & v0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p23_hpc22_G4_mul1_G16_mul0_G256_inv0 = (u1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p3_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p23_hpc22_G4_mul1_G16_mul0_G256_inv0);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q1_G4_mul1_G16_mul0_G256_inv0 = (q1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign z4025_assgn4025 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul0_G256_inv0 = (p1_G4_mul1_G16_mul0_G256_inv0 << z899_assgn899);
    assign z4029_assgn4029 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << z901_assgn901);
    assign p0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul1_G16_mul0_G256_inv0 | q1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p1_G16_mul0_G256_inv0 = (p1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign r00_G4_mul2_G16_mul0_G256_inv0 = (r60_G16_mul0_G256_inv0 % z3_assgn3);
    assign r10_G4_mul2_G16_mul0_G256_inv0 = (r70_G16_mul0_G256_inv0 % z3_assgn3);
    assign r20_G4_mul2_G16_mul0_G256_inv0 = (r80_G16_mul0_G256_inv0 % z3_assgn3);
    assign z4047_assgn4047 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & z917_assgn917);
    assign z4051_assgn4051 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & z919_assgn919);
    assign z4055_assgn4055 = dec_1_inp;
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> z921_assgn921);
    assign z4059_assgn4059 = dec_1_inp;
    assign a1_G4_mul2_G16_mul0_G256_inv0 = (a1_0_G4_mul2_G16_mul0_G256_inv0 >> z923_assgn923);
    assign z4063_assgn4063 = dec_1_inp;
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & z925_assgn925);
    assign z4067_assgn4067 = dec_1_inp;
    assign b1_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & z927_assgn927);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul0_G256_inv0 = (c1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0_reg ^ d0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign axorb_1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ b1_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0_reg ^ d1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign r0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0 = !axorb_0_G4_mul2_G16_mul0_G256_inv0;
    assign a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0 = !axorb_1_G4_mul2_G16_mul0_G256_inv0;
    assign z4097_assgn4097 = r0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    assign u0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0 & z955_assgn955);
    assign z4101_assgn4101 = r0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    assign u1_hpc20_G4_mul2_G16_mul0_G256_inv0 = (a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0 & z957_assgn957);
    assign v0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (cxord_0_G4_mul2_G16_mul0_G256_inv0_reg ^ r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign v1_hpc20_G4_mul2_G16_mul0_G256_inv0 = (cxord_1_G4_mul2_G16_mul0_G256_inv0_reg ^ r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign z4109_assgn4109 = cxord_0_G4_mul2_G16_mul0_G256_inv0;
    assign p0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 & z963_assgn963);
    assign p1_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 & v1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p01_hpc20_G4_mul2_G16_mul0_G256_inv0 = (u0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul0_G256_inv0 = (p0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p01_hpc20_G4_mul2_G16_mul0_G256_inv0);
    assign z4119_assgn4119 = cxord_1_G4_mul2_G16_mul0_G256_inv0;
    assign p2_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0 & z971_assgn971);
    assign p3_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0 & v0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p23_hpc20_G4_mul2_G16_mul0_G256_inv0 = (u1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p3_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p23_hpc20_G4_mul2_G16_mul0_G256_inv0);
    assign r0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0 = !a0_G4_mul2_G16_mul0_G256_inv0;
    assign a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0 = !a1_G4_mul2_G16_mul0_G256_inv0;
    assign z4135_assgn4135 = r0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    assign u0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0 & z985_assgn985);
    assign z4139_assgn4139 = r0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    assign u1_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0 & z987_assgn987);
    assign z4143_assgn4143 = c0_G4_mul2_G16_mul0_G256_inv0;
    assign v0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (z990_assgn990 ^ r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign z4147_assgn4147 = c1_G4_mul2_G16_mul0_G256_inv0;
    assign v1_hpc21_G4_mul2_G16_mul0_G256_inv0 = (z992_assgn992 ^ r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign z4151_assgn4151 = c0_G4_mul2_G16_mul0_G256_inv0;
    assign p0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 & z993_assgn993);
    assign p1_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 & v1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p01_hpc21_G4_mul2_G16_mul0_G256_inv0 = (u0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (p0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p01_hpc21_G4_mul2_G16_mul0_G256_inv0);
    assign z4161_assgn4161 = c1_G4_mul2_G16_mul0_G256_inv0;
    assign p2_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 & z1001_assgn1001);
    assign p3_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 & v0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p23_hpc21_G4_mul2_G16_mul0_G256_inv0 = (u1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p3_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p23_hpc21_G4_mul2_G16_mul0_G256_inv0);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_G4_mul2_G16_mul0_G256_inv0 = (p1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign r0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp_reg);
    assign a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0 = !b0_G4_mul2_G16_mul0_G256_inv0;
    assign a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0 = !b1_G4_mul2_G16_mul0_G256_inv0;
    assign z4181_assgn4181 = r0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    assign u0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0 & z1019_assgn1019);
    assign z4185_assgn4185 = r0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    assign u1_hpc22_G4_mul2_G16_mul0_G256_inv0 = (a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0 & z1021_assgn1021);
    assign z4189_assgn4189 = d0_G4_mul2_G16_mul0_G256_inv0;
    assign v0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (z1024_assgn1024 ^ r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign z4193_assgn4193 = d1_G4_mul2_G16_mul0_G256_inv0;
    assign v1_hpc22_G4_mul2_G16_mul0_G256_inv0 = (z1026_assgn1026 ^ r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign z4197_assgn4197 = d0_G4_mul2_G16_mul0_G256_inv0;
    assign p0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 & z1027_assgn1027);
    assign p1_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 & v1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p01_hpc22_G4_mul2_G16_mul0_G256_inv0 = (u0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (p0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p01_hpc22_G4_mul2_G16_mul0_G256_inv0);
    assign z4207_assgn4207 = d1_G4_mul2_G16_mul0_G256_inv0;
    assign p2_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0 & z1035_assgn1035);
    assign p3_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0 & v0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p23_hpc22_G4_mul2_G16_mul0_G256_inv0 = (u1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p3_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p23_hpc22_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q1_G4_mul2_G16_mul0_G256_inv0 = (q1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign z4221_assgn4221 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul0_G256_inv0 = (p1_G4_mul2_G16_mul0_G256_inv0 << z1047_assgn1047);
    assign z4225_assgn4225 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << z1049_assgn1049);
    assign q0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul2_G16_mul0_G256_inv0 | q1_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign q1_G16_mul0_G256_inv0 = (q1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign z4237_assgn4237 = dec_2_inp;
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << z1059_assgn1059);
    assign z4241_assgn4241 = dec_2_inp;
    assign p1ls2_G16_mul0_G256_inv0 = (p1_G16_mul0_G256_inv0 << z1061_assgn1061);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign d1_G256_inv0 = (p1ls2_G16_mul0_G256_inv0 | q1_G16_mul0_G256_inv0);
    assign c0xord0_G256_inv0 = (c0_G256_inv0 ^ d0_G256_inv0);
    assign c1xord1_G256_inv0 = (c1_G256_inv0 ^ d1_G256_inv0);
    assign z4253_assgn4253 = z1_assgn1;
    assign r00_G16_inv0_G256_inv0 = (r9_inp % z1071_assgn1071);
    assign z4257_assgn4257 = z1_assgn1;
    assign r10_G16_inv0_G256_inv0 = (r10_inp % z1073_assgn1073);
    assign z4261_assgn4261 = z1_assgn1;
    assign r20_G16_inv0_G256_inv0 = (r11_inp % z1075_assgn1075);
    assign z4265_assgn4265 = z1_assgn1;
    assign r30_G16_inv0_G256_inv0 = (r12_inp % z1077_assgn1077);
    assign z4269_assgn4269 = z1_assgn1;
    assign r40_G16_inv0_G256_inv0 = (r13_inp % z1079_assgn1079);
    assign z4273_assgn4273 = z1_assgn1;
    assign r50_G16_inv0_G256_inv0 = (r14_inp % z1081_assgn1081);
    assign z4277_assgn4277 = z1_assgn1;
    assign r60_G16_inv0_G256_inv0 = (r15_inp % z1083_assgn1083);
    assign z4281_assgn4281 = z1_assgn1;
    assign r70_G16_inv0_G256_inv0 = (r16_inp % z1085_assgn1085);
    assign z4285_assgn4285 = z1_assgn1;
    assign r80_G16_inv0_G256_inv0 = (r17_inp % z1087_assgn1087);
    assign z4289_assgn4289 = dec_12_inp;
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0_reg & z1089_assgn1089);
    assign z4293_assgn4293 = dec_12_inp;
    assign a1_0_G16_inv0_G256_inv0 = (c1xord1_G256_inv0_reg & z1091_assgn1091);
    assign z4297_assgn4297 = dec_2_inp;
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> z1093_assgn1093);
    assign z4301_assgn4301 = dec_2_inp;
    assign a1_G16_inv0_G256_inv0 = (a1_0_G16_inv0_G256_inv0 >> z1095_assgn1095);
    assign z4305_assgn4305 = dec_3_inp;
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & z1097_assgn1097);
    assign z4309_assgn4309 = dec_3_inp;
    assign b1_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1099_assgn1099);
    assign z4313_assgn4313 = b0_G16_inv0_G256_inv0;
    assign z4315_assgn4315 = a0_G16_inv0_G256_inv0;
    assign a0xorb0_G16_inv0_G256_inv0 = (z1102_assgn1102 ^ z1101_assgn1101);
    assign z4319_assgn4319 = b1_G16_inv0_G256_inv0;
    assign z4321_assgn4321 = a1_G16_inv0_G256_inv0;
    assign a1xorb1_G16_inv0_G256_inv0 = (z1104_assgn1104 ^ z1103_assgn1103);
    assign z4325_assgn4325 = dec_2_inp;
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & z1105_assgn1105);
    assign z4329_assgn4329 = dec_2_inp;
    assign a1_0_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1107_assgn1107);
    assign z4333_assgn4333 = dec_1_inp;
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> z1109_assgn1109);
    assign z4337_assgn4337 = dec_1_inp;
    assign a1_G4_sq2_G16_inv0_G256_inv0 = (a1_0_G4_sq2_G16_inv0_G256_inv0 >> z1111_assgn1111);
    assign z4341_assgn4341 = dec_1_inp;
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & z1113_assgn1113);
    assign z4345_assgn4345 = dec_1_inp;
    assign b1_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1115_assgn1115);
    assign z4349_assgn4349 = dec_1_inp;
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << z1117_assgn1117);
    assign z4353_assgn4353 = dec_1_inp;
    assign b1ls1_G4_sq2_G16_inv0_G256_inv0 = (b1_G4_sq2_G16_inv0_G256_inv0 << z1119_assgn1119);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign c1_0_G16_inv0_G256_inv0 = (b1ls1_G4_sq2_G16_inv0_G256_inv0 | a1_G4_sq2_G16_inv0_G256_inv0);
    assign z4361_assgn4361 = dec_2_inp;
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & z1125_assgn1125);
    assign z4365_assgn4365 = dec_2_inp;
    assign a1_0_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1127_assgn1127);
    assign z4369_assgn4369 = dec_1_inp;
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1129_assgn1129);
    assign z4373_assgn4373 = dec_1_inp;
    assign a1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1131_assgn1131);
    assign z4377_assgn4377 = dec_1_inp;
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & z1133_assgn1133);
    assign z4381_assgn4381 = dec_1_inp;
    assign b1_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1135_assgn1135);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign p1_G4_scl_N1_G16_inv0_G256_inv0 = b1_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign q1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_G4_scl_N1_G16_inv0_G256_inv0 ^ b1_G4_scl_N1_G16_inv0_G256_inv0);
    assign z4393_assgn4393 = dec_1_inp;
    assign p1ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p1_G4_scl_N1_G16_inv0_G256_inv0 << z1145_assgn1145);
    assign z4397_assgn4397 = dec_1_inp;
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << z1147_assgn1147);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign c1_G16_inv0_G256_inv0 = (p1ls1_G4_scl_N1_G16_inv0_G256_inv0 | q1_G4_scl_N1_G16_inv0_G256_inv0);
    assign z4405_assgn4405 = z3_assgn3;
    assign r00_G4_mul3_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % z1153_assgn1153);
    assign z4409_assgn4409 = z3_assgn3;
    assign r10_G4_mul3_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % z1155_assgn1155);
    assign z4413_assgn4413 = z3_assgn3;
    assign r20_G4_mul3_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % z1157_assgn1157);
    assign z4417_assgn4417 = dec_2_inp;
    assign z4419_assgn4419 = a0_G16_inv0_G256_inv0;
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (z1160_assgn1160 & z1159_assgn1159);
    assign z4423_assgn4423 = dec_2_inp;
    assign z4425_assgn4425 = a1_G16_inv0_G256_inv0;
    assign a1_0_G4_mul3_G16_inv0_G256_inv0 = (z1162_assgn1162 & z1161_assgn1161);
    assign z4429_assgn4429 = dec_1_inp;
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> z1163_assgn1163);
    assign z4433_assgn4433 = dec_1_inp;
    assign a1_G4_mul3_G16_inv0_G256_inv0 = (a1_0_G4_mul3_G16_inv0_G256_inv0 >> z1165_assgn1165);
    assign z4437_assgn4437 = dec_1_inp;
    assign z4439_assgn4439 = a0_G16_inv0_G256_inv0;
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (z1168_assgn1168 & z1167_assgn1167);
    assign z4443_assgn4443 = dec_1_inp;
    assign z4445_assgn4445 = a1_G16_inv0_G256_inv0;
    assign b1_G4_mul3_G16_inv0_G256_inv0 = (z1170_assgn1170 & z1169_assgn1169);
    assign z4449_assgn4449 = dec_2_inp;
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1171_assgn1171);
    assign z4453_assgn4453 = dec_2_inp;
    assign c1_0_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1173_assgn1173);
    assign z4457_assgn4457 = dec_1_inp;
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> z1175_assgn1175);
    assign z4461_assgn4461 = dec_1_inp;
    assign c1_G4_mul3_G16_inv0_G256_inv0 = (c1_0_G4_mul3_G16_inv0_G256_inv0 >> z1177_assgn1177);
    assign z4465_assgn4465 = dec_1_inp;
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1179_assgn1179);
    assign z4469_assgn4469 = dec_1_inp;
    assign d1_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1181_assgn1181);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0_reg ^ d0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign axorb_1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ b1_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0_reg ^ d1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4481_assgn4481 = dec_2_inp;
    assign r0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % z1191_assgn1191);
    assign a0_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 = !axorb_0_G4_mul3_G16_inv0_G256_inv0;
    assign a1_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 = !axorb_1_G4_mul3_G16_inv0_G256_inv0;
    assign z4489_assgn4489 = r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign u0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (a0_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 & z1197_assgn1197);
    assign z4493_assgn4493 = r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign u1_hpc20_G4_mul3_G16_inv0_G256_inv0 = (a1_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 & z1199_assgn1199);
    assign v0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (cxord_0_G4_mul3_G16_inv0_G256_inv0_reg ^ r0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign v1_hpc20_G4_mul3_G16_inv0_G256_inv0 = (cxord_1_G4_mul3_G16_inv0_G256_inv0_reg ^ r0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4501_assgn4501 = cxord_0_G4_mul3_G16_inv0_G256_inv0;
    assign p0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 & z1205_assgn1205);
    assign p1_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 & v1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p01_hpc20_G4_mul3_G16_inv0_G256_inv0 = (u0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul3_G16_inv0_G256_inv0 = (p0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg ^ p01_hpc20_G4_mul3_G16_inv0_G256_inv0);
    assign z4511_assgn4511 = cxord_1_G4_mul3_G16_inv0_G256_inv0;
    assign p2_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0 & z1213_assgn1213);
    assign p3_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0 & v0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p23_hpc20_G4_mul3_G16_inv0_G256_inv0 = (u1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg ^ p3_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc20_G4_mul3_G16_inv0_G256_inv0_reg ^ p23_hpc20_G4_mul3_G16_inv0_G256_inv0);
    assign z4521_assgn4521 = dec_2_inp;
    assign r0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % z1221_assgn1221);
    assign a0_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 = !a0_G4_mul3_G16_inv0_G256_inv0;
    assign a1_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 = !a1_G4_mul3_G16_inv0_G256_inv0;
    assign z4529_assgn4529 = r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign u0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a0_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 & z1227_assgn1227);
    assign z4533_assgn4533 = r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign u1_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a1_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 & z1229_assgn1229);
    assign z4537_assgn4537 = c0_G4_mul3_G16_inv0_G256_inv0;
    assign v0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (z1232_assgn1232 ^ r0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4541_assgn4541 = c1_G4_mul3_G16_inv0_G256_inv0;
    assign v1_hpc21_G4_mul3_G16_inv0_G256_inv0 = (z1234_assgn1234 ^ r0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4545_assgn4545 = c0_G4_mul3_G16_inv0_G256_inv0;
    assign p0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 & z1235_assgn1235);
    assign p1_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 & v1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p01_hpc21_G4_mul3_G16_inv0_G256_inv0 = (u0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (p0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg ^ p01_hpc21_G4_mul3_G16_inv0_G256_inv0);
    assign z4555_assgn4555 = c1_G4_mul3_G16_inv0_G256_inv0;
    assign p2_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 & z1243_assgn1243);
    assign p3_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 & v0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p23_hpc21_G4_mul3_G16_inv0_G256_inv0 = (u1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg ^ p3_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc21_G4_mul3_G16_inv0_G256_inv0_reg ^ p23_hpc21_G4_mul3_G16_inv0_G256_inv0);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_G4_mul3_G16_inv0_G256_inv0 = (p1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign z4569_assgn4569 = dec_2_inp;
    assign r0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % z1255_assgn1255);
    assign a0_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 = !b0_G4_mul3_G16_inv0_G256_inv0;
    assign a1_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 = !b1_G4_mul3_G16_inv0_G256_inv0;
    assign z4577_assgn4577 = r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign u0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (a0_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 & z1261_assgn1261);
    assign z4581_assgn4581 = r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign u1_hpc22_G4_mul3_G16_inv0_G256_inv0 = (a1_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 & z1263_assgn1263);
    assign z4585_assgn4585 = d0_G4_mul3_G16_inv0_G256_inv0;
    assign v0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (z1266_assgn1266 ^ r0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4589_assgn4589 = d1_G4_mul3_G16_inv0_G256_inv0;
    assign v1_hpc22_G4_mul3_G16_inv0_G256_inv0 = (z1268_assgn1268 ^ r0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4593_assgn4593 = d0_G4_mul3_G16_inv0_G256_inv0;
    assign p0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 & z1269_assgn1269);
    assign p1_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 & v1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p01_hpc22_G4_mul3_G16_inv0_G256_inv0 = (u0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (p0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg ^ p01_hpc22_G4_mul3_G16_inv0_G256_inv0);
    assign z4603_assgn4603 = d1_G4_mul3_G16_inv0_G256_inv0;
    assign p2_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0 & z1277_assgn1277);
    assign p3_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0 & v0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p23_hpc22_G4_mul3_G16_inv0_G256_inv0 = (u1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg ^ p3_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc22_G4_mul3_G16_inv0_G256_inv0_reg ^ p23_hpc22_G4_mul3_G16_inv0_G256_inv0);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q1_G4_mul3_G16_inv0_G256_inv0 = (q1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign z4617_assgn4617 = dec_1_inp;
    assign p1ls1_G4_mul3_G16_inv0_G256_inv0 = (p1_G4_mul3_G16_inv0_G256_inv0 << z1289_assgn1289);
    assign z4621_assgn4621 = dec_1_inp;
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << z1291_assgn1291);
    assign d0_G16_inv0_G256_inv0 = (p1ls1_G4_mul3_G16_inv0_G256_inv0 | q1_G4_mul3_G16_inv0_G256_inv0);
    assign d1_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign c0xord0_G16_inv0_G256_inv0 = (c0_G16_inv0_G256_inv0 ^ d0_G16_inv0_G256_inv0);
    assign c1xord1_G16_inv0_G256_inv0 = (c1_G16_inv0_G256_inv0 ^ d1_G16_inv0_G256_inv0);
    assign z4633_assgn4633 = dec_2_inp;
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1301_assgn1301);
    assign z4637_assgn4637 = dec_2_inp;
    assign a1_0_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1303_assgn1303);
    assign z4641_assgn4641 = dec_1_inp;
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> z1305_assgn1305);
    assign z4645_assgn4645 = dec_1_inp;
    assign a1_G4_sq3_G16_inv0_G256_inv0 = (a1_0_G4_sq3_G16_inv0_G256_inv0 >> z1307_assgn1307);
    assign z4649_assgn4649 = dec_1_inp;
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1309_assgn1309);
    assign z4653_assgn4653 = dec_1_inp;
    assign b1_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1311_assgn1311);
    assign z4657_assgn4657 = dec_1_inp;
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << z1313_assgn1313);
    assign z4661_assgn4661 = dec_1_inp;
    assign b1ls1_G4_sq3_G16_inv0_G256_inv0 = (b1_G4_sq3_G16_inv0_G256_inv0 << z1315_assgn1315);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign e1_G16_inv0_G256_inv0 = (b1ls1_G4_sq3_G16_inv0_G256_inv0 | a1_G4_sq3_G16_inv0_G256_inv0);
    assign z4669_assgn4669 = z3_assgn3;
    assign r00_G4_mul4_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % z1321_assgn1321);
    assign z4673_assgn4673 = z3_assgn3;
    assign r10_G4_mul4_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % z1323_assgn1323);
    assign z4677_assgn4677 = z3_assgn3;
    assign r20_G4_mul4_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % z1325_assgn1325);
    assign z4681_assgn4681 = dec_2_inp;
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1327_assgn1327);
    assign z4685_assgn4685 = dec_2_inp;
    assign a1_0_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1329_assgn1329);
    assign z4689_assgn4689 = dec_1_inp;
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> z1331_assgn1331);
    assign z4693_assgn4693 = dec_1_inp;
    assign a1_G4_mul4_G16_inv0_G256_inv0 = (a1_0_G4_mul4_G16_inv0_G256_inv0 >> z1333_assgn1333);
    assign z4697_assgn4697 = dec_1_inp;
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1335_assgn1335);
    assign z4701_assgn4701 = dec_1_inp;
    assign b1_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1337_assgn1337);
    assign z4705_assgn4705 = dec_2_inp;
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0_reg & z1339_assgn1339);
    assign z4709_assgn4709 = dec_2_inp;
    assign c1_0_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0_reg & z1341_assgn1341);
    assign z4713_assgn4713 = dec_1_inp;
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> z1343_assgn1343);
    assign z4717_assgn4717 = dec_1_inp;
    assign c1_G4_mul4_G16_inv0_G256_inv0 = (c1_0_G4_mul4_G16_inv0_G256_inv0 >> z1345_assgn1345);
    assign z4721_assgn4721 = dec_1_inp;
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0_reg & z1347_assgn1347);
    assign z4725_assgn4725 = dec_1_inp;
    assign d1_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0_reg & z1349_assgn1349);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0_reg ^ d0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign axorb_1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ b1_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0_reg ^ d1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z4737_assgn4737 = dec_2_inp;
    assign r0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % z1359_assgn1359);
    assign a0_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 = !axorb_0_G4_mul4_G16_inv0_G256_inv0;
    assign a1_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 = !axorb_1_G4_mul4_G16_inv0_G256_inv0;
    assign z4745_assgn4745 = r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign u0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (a0_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 & z1365_assgn1365);
    assign z4749_assgn4749 = r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign u1_hpc20_G4_mul4_G16_inv0_G256_inv0 = (a1_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 & z1367_assgn1367);
    assign v0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (cxord_0_G4_mul4_G16_inv0_G256_inv0_reg ^ r0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign v1_hpc20_G4_mul4_G16_inv0_G256_inv0 = (cxord_1_G4_mul4_G16_inv0_G256_inv0_reg ^ r0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z4757_assgn4757 = cxord_0_G4_mul4_G16_inv0_G256_inv0;
    assign p0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & z1373_assgn1373);
    assign p1_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & v1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p01_hpc20_G4_mul4_G16_inv0_G256_inv0 = (u0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul4_G16_inv0_G256_inv0 = (p0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p01_hpc20_G4_mul4_G16_inv0_G256_inv0);
    assign z4767_assgn4767 = cxord_1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & z1381_assgn1381);
    assign p3_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & v0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p23_hpc20_G4_mul4_G16_inv0_G256_inv0 = (u1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p3_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p23_hpc20_G4_mul4_G16_inv0_G256_inv0);
    assign z4777_assgn4777 = dec_2_inp;
    assign r0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % z1389_assgn1389);
    assign a0_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 = !a0_G4_mul4_G16_inv0_G256_inv0;
    assign a1_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 = !a1_G4_mul4_G16_inv0_G256_inv0;
    assign z4785_assgn4785 = r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign u0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a0_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 & z1395_assgn1395);
    assign z4789_assgn4789 = r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign u1_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a1_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 & z1397_assgn1397);
    assign z4793_assgn4793 = c0_G4_mul4_G16_inv0_G256_inv0;
    assign v0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (z1400_assgn1400 ^ r0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z4797_assgn4797 = c1_G4_mul4_G16_inv0_G256_inv0;
    assign v1_hpc21_G4_mul4_G16_inv0_G256_inv0 = (z1402_assgn1402 ^ r0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z4801_assgn4801 = c0_G4_mul4_G16_inv0_G256_inv0;
    assign p0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & z1403_assgn1403);
    assign p1_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & v1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p01_hpc21_G4_mul4_G16_inv0_G256_inv0 = (u0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (p0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p01_hpc21_G4_mul4_G16_inv0_G256_inv0);
    assign z4811_assgn4811 = c1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & z1411_assgn1411);
    assign p3_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & v0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p23_hpc21_G4_mul4_G16_inv0_G256_inv0 = (u1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p3_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p23_hpc21_G4_mul4_G16_inv0_G256_inv0);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G4_mul4_G16_inv0_G256_inv0 = (p1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign z4825_assgn4825 = dec_2_inp;
    assign r0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % z1423_assgn1423);
    assign a0_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 = !b0_G4_mul4_G16_inv0_G256_inv0;
    assign a1_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 = !b1_G4_mul4_G16_inv0_G256_inv0;
    assign z4833_assgn4833 = r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign u0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (a0_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 & z1429_assgn1429);
    assign z4837_assgn4837 = r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign u1_hpc22_G4_mul4_G16_inv0_G256_inv0 = (a1_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 & z1431_assgn1431);
    assign z4841_assgn4841 = d0_G4_mul4_G16_inv0_G256_inv0;
    assign v0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (z1434_assgn1434 ^ r0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z4845_assgn4845 = d1_G4_mul4_G16_inv0_G256_inv0;
    assign v1_hpc22_G4_mul4_G16_inv0_G256_inv0 = (z1436_assgn1436 ^ r0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z4849_assgn4849 = d0_G4_mul4_G16_inv0_G256_inv0;
    assign p0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & z1437_assgn1437);
    assign p1_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & v1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p01_hpc22_G4_mul4_G16_inv0_G256_inv0 = (u0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (p0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p01_hpc22_G4_mul4_G16_inv0_G256_inv0);
    assign z4859_assgn4859 = d1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & z1445_assgn1445);
    assign p3_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & v0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p23_hpc22_G4_mul4_G16_inv0_G256_inv0 = (u1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p3_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p23_hpc22_G4_mul4_G16_inv0_G256_inv0);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q1_G4_mul4_G16_inv0_G256_inv0 = (q1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign z4873_assgn4873 = dec_1_inp;
    assign p1ls1_G4_mul4_G16_inv0_G256_inv0 = (p1_G4_mul4_G16_inv0_G256_inv0 << z1457_assgn1457);
    assign z4877_assgn4877 = dec_1_inp;
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << z1459_assgn1459);
    assign p0_G16_inv0_G256_inv0 = (p1ls1_G4_mul4_G16_inv0_G256_inv0 | q1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign z4885_assgn4885 = z3_assgn3;
    assign r00_G4_mul5_G16_inv0_G256_inv0 = (r60_G16_inv0_G256_inv0 % z1465_assgn1465);
    assign z4889_assgn4889 = z3_assgn3;
    assign r10_G4_mul5_G16_inv0_G256_inv0 = (r70_G16_inv0_G256_inv0 % z1467_assgn1467);
    assign z4893_assgn4893 = z3_assgn3;
    assign r20_G4_mul5_G16_inv0_G256_inv0 = (r80_G16_inv0_G256_inv0 % z1469_assgn1469);
    assign z4897_assgn4897 = dec_2_inp;
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1471_assgn1471);
    assign z4901_assgn4901 = dec_2_inp;
    assign a1_0_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1473_assgn1473);
    assign z4905_assgn4905 = dec_1_inp;
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> z1475_assgn1475);
    assign z4909_assgn4909 = dec_1_inp;
    assign a1_G4_mul5_G16_inv0_G256_inv0 = (a1_0_G4_mul5_G16_inv0_G256_inv0 >> z1477_assgn1477);
    assign z4913_assgn4913 = dec_1_inp;
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1479_assgn1479);
    assign z4917_assgn4917 = dec_1_inp;
    assign b1_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1481_assgn1481);
    assign z4921_assgn4921 = dec_2_inp;
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1483_assgn1483);
    assign z4925_assgn4925 = dec_2_inp;
    assign c1_0_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1485_assgn1485);
    assign z4929_assgn4929 = dec_1_inp;
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> z1487_assgn1487);
    assign z4933_assgn4933 = dec_1_inp;
    assign c1_G4_mul5_G16_inv0_G256_inv0 = (c1_0_G4_mul5_G16_inv0_G256_inv0 >> z1489_assgn1489);
    assign z4937_assgn4937 = dec_1_inp;
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1491_assgn1491);
    assign z4941_assgn4941 = dec_1_inp;
    assign d1_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1493_assgn1493);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0_reg ^ d0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign axorb_1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ b1_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0_reg ^ d1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z4953_assgn4953 = dec_2_inp;
    assign r0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % z1503_assgn1503);
    assign a0_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 = !axorb_0_G4_mul5_G16_inv0_G256_inv0;
    assign a1_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 = !axorb_1_G4_mul5_G16_inv0_G256_inv0;
    assign z4961_assgn4961 = r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign u0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (a0_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 & z1509_assgn1509);
    assign z4965_assgn4965 = r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign u1_hpc20_G4_mul5_G16_inv0_G256_inv0 = (a1_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 & z1511_assgn1511);
    assign v0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (cxord_0_G4_mul5_G16_inv0_G256_inv0_reg ^ r0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign v1_hpc20_G4_mul5_G16_inv0_G256_inv0 = (cxord_1_G4_mul5_G16_inv0_G256_inv0_reg ^ r0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z4973_assgn4973 = cxord_0_G4_mul5_G16_inv0_G256_inv0;
    assign p0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & z1517_assgn1517);
    assign p1_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & v1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p01_hpc20_G4_mul5_G16_inv0_G256_inv0 = (u0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul5_G16_inv0_G256_inv0 = (p0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p01_hpc20_G4_mul5_G16_inv0_G256_inv0);
    assign z4983_assgn4983 = cxord_1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & z1525_assgn1525);
    assign p3_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & v0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p23_hpc20_G4_mul5_G16_inv0_G256_inv0 = (u1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p3_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p23_hpc20_G4_mul5_G16_inv0_G256_inv0);
    assign z4993_assgn4993 = dec_2_inp;
    assign r0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % z1533_assgn1533);
    assign a0_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 = !a0_G4_mul5_G16_inv0_G256_inv0;
    assign a1_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 = !a1_G4_mul5_G16_inv0_G256_inv0;
    assign z5001_assgn5001 = r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign u0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a0_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 & z1539_assgn1539);
    assign z5005_assgn5005 = r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign u1_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a1_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 & z1541_assgn1541);
    assign z5009_assgn5009 = c0_G4_mul5_G16_inv0_G256_inv0;
    assign v0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (z1544_assgn1544 ^ r0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5013_assgn5013 = c1_G4_mul5_G16_inv0_G256_inv0;
    assign v1_hpc21_G4_mul5_G16_inv0_G256_inv0 = (z1546_assgn1546 ^ r0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5017_assgn5017 = c0_G4_mul5_G16_inv0_G256_inv0;
    assign p0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & z1547_assgn1547);
    assign p1_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & v1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p01_hpc21_G4_mul5_G16_inv0_G256_inv0 = (u0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (p0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p01_hpc21_G4_mul5_G16_inv0_G256_inv0);
    assign z5027_assgn5027 = c1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & z1555_assgn1555);
    assign p3_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & v0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p23_hpc21_G4_mul5_G16_inv0_G256_inv0 = (u1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p3_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p23_hpc21_G4_mul5_G16_inv0_G256_inv0);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_G4_mul5_G16_inv0_G256_inv0 = (p1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign z5041_assgn5041 = dec_2_inp;
    assign r0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % z1567_assgn1567);
    assign a0_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 = !b0_G4_mul5_G16_inv0_G256_inv0;
    assign a1_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 = !b1_G4_mul5_G16_inv0_G256_inv0;
    assign z5049_assgn5049 = r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign u0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (a0_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 & z1573_assgn1573);
    assign z5053_assgn5053 = r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign u1_hpc22_G4_mul5_G16_inv0_G256_inv0 = (a1_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 & z1575_assgn1575);
    assign z5057_assgn5057 = d0_G4_mul5_G16_inv0_G256_inv0;
    assign v0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (z1578_assgn1578 ^ r0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5061_assgn5061 = d1_G4_mul5_G16_inv0_G256_inv0;
    assign v1_hpc22_G4_mul5_G16_inv0_G256_inv0 = (z1580_assgn1580 ^ r0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5065_assgn5065 = d0_G4_mul5_G16_inv0_G256_inv0;
    assign p0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & z1581_assgn1581);
    assign p1_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & v1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p01_hpc22_G4_mul5_G16_inv0_G256_inv0 = (u0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (p0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p01_hpc22_G4_mul5_G16_inv0_G256_inv0);
    assign z5075_assgn5075 = d1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & z1589_assgn1589);
    assign p3_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & v0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p23_hpc22_G4_mul5_G16_inv0_G256_inv0 = (u1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p3_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p23_hpc22_G4_mul5_G16_inv0_G256_inv0);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G4_mul5_G16_inv0_G256_inv0 = (q1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign z5089_assgn5089 = dec_1_inp;
    assign p1ls1_G4_mul5_G16_inv0_G256_inv0 = (p1_G4_mul5_G16_inv0_G256_inv0 << z1601_assgn1601);
    assign z5093_assgn5093 = dec_1_inp;
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << z1603_assgn1603);
    assign q0_G16_inv0_G256_inv0 = (p1ls1_G4_mul5_G16_inv0_G256_inv0 | q1_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign z5101_assgn5101 = dec_2_inp;
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << z1609_assgn1609);
    assign z5105_assgn5105 = dec_2_inp;
    assign p1ls2_G16_inv0_G256_inv0 = (p1_G16_inv0_G256_inv0 << z1611_assgn1611);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign e1_G256_inv0 = (p1ls2_G16_inv0_G256_inv0 | q1_G16_inv0_G256_inv0);
    assign z5113_assgn5113 = z1_assgn1;
    assign r00_G16_mul1_G256_inv0 = (r18_inp % z1617_assgn1617);
    assign z5117_assgn5117 = z1_assgn1;
    assign r10_G16_mul1_G256_inv0 = (r19_inp % z1619_assgn1619);
    assign z5121_assgn5121 = z1_assgn1;
    assign r20_G16_mul1_G256_inv0 = (r20_inp % z1621_assgn1621);
    assign z5125_assgn5125 = z1_assgn1;
    assign r30_G16_mul1_G256_inv0 = (r21_inp % z1623_assgn1623);
    assign z5129_assgn5129 = z1_assgn1;
    assign r40_G16_mul1_G256_inv0 = (r22_inp % z1625_assgn1625);
    assign z5133_assgn5133 = z1_assgn1;
    assign r50_G16_mul1_G256_inv0 = (r23_inp % z1627_assgn1627);
    assign z5137_assgn5137 = z1_assgn1;
    assign r60_G16_mul1_G256_inv0 = (r24_inp % z1629_assgn1629);
    assign z5141_assgn5141 = z1_assgn1;
    assign r70_G16_mul1_G256_inv0 = (r25_inp % z1631_assgn1631);
    assign z5145_assgn5145 = z1_assgn1;
    assign r80_G16_mul1_G256_inv0 = (r26_inp % z1633_assgn1633);
    assign z5149_assgn5149 = dec_12_inp;
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1635_assgn1635);
    assign z5153_assgn5153 = dec_12_inp;
    assign a1_0_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1637_assgn1637);
    assign z5157_assgn5157 = dec_2_inp;
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> z1639_assgn1639);
    assign z5161_assgn5161 = dec_2_inp;
    assign a1_G16_mul1_G256_inv0 = (a1_0_G16_mul1_G256_inv0 >> z1641_assgn1641);
    assign z5165_assgn5165 = dec_3_inp;
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1643_assgn1643);
    assign z5169_assgn5169 = dec_3_inp;
    assign b1_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1645_assgn1645);
    assign z5173_assgn5173 = dec_12_inp;
    assign z5175_assgn5175 = b0_G256_inv0;
    assign c0_0_G16_mul1_G256_inv0 = (z1648_assgn1648 & z1647_assgn1647);
    assign z5179_assgn5179 = dec_12_inp;
    assign z5181_assgn5181 = b1_G256_inv0;
    assign c1_0_G16_mul1_G256_inv0 = (z1650_assgn1650 & z1649_assgn1649);
    assign z5185_assgn5185 = dec_2_inp;
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> z1651_assgn1651);
    assign z5189_assgn5189 = dec_2_inp;
    assign c1_G16_mul1_G256_inv0 = (c1_0_G16_mul1_G256_inv0 >> z1653_assgn1653);
    assign z5193_assgn5193 = dec_3_inp;
    assign z5195_assgn5195 = b0_G256_inv0;
    assign d0_G16_mul1_G256_inv0 = (z1656_assgn1656 & z1655_assgn1655);
    assign z5199_assgn5199 = dec_3_inp;
    assign z5201_assgn5201 = b1_G256_inv0;
    assign d1_G16_mul1_G256_inv0 = (z1658_assgn1658 & z1657_assgn1657);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign axorb_1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 ^ b1_G16_mul1_G256_inv0);
    assign cxord_1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 ^ d1_G16_mul1_G256_inv0);
    assign z5213_assgn5213 = z3_assgn3;
    assign r00_G4_mul0_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % z1667_assgn1667);
    assign z5217_assgn5217 = z3_assgn3;
    assign r10_G4_mul0_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % z1669_assgn1669);
    assign z5221_assgn5221 = z3_assgn3;
    assign r20_G4_mul0_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % z1671_assgn1671);
    assign z5225_assgn5225 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1673_assgn1673);
    assign z5229_assgn5229 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1675_assgn1675);
    assign z5233_assgn5233 = dec_1_inp;
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> z1677_assgn1677);
    assign z5237_assgn5237 = dec_1_inp;
    assign a1_G4_mul0_G16_mul1_G256_inv0 = (a1_0_G4_mul0_G16_mul1_G256_inv0 >> z1679_assgn1679);
    assign z5241_assgn5241 = dec_1_inp;
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1681_assgn1681);
    assign z5245_assgn5245 = dec_1_inp;
    assign b1_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1683_assgn1683);
    assign z5249_assgn5249 = dec_2_inp;
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & z1685_assgn1685);
    assign z5253_assgn5253 = dec_2_inp;
    assign c1_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & z1687_assgn1687);
    assign z5257_assgn5257 = dec_1_inp;
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> z1689_assgn1689);
    assign z5261_assgn5261 = dec_1_inp;
    assign c1_G4_mul0_G16_mul1_G256_inv0 = (c1_0_G4_mul0_G16_mul1_G256_inv0 >> z1691_assgn1691);
    assign z5265_assgn5265 = dec_1_inp;
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & z1693_assgn1693);
    assign z5269_assgn5269 = dec_1_inp;
    assign d1_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & z1695_assgn1695);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0_reg ^ d0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign axorb_1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ b1_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0_reg ^ d1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5281_assgn5281 = dec_2_inp;
    assign r0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % z1705_assgn1705);
    assign a0_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 = !axorb_0_G4_mul0_G16_mul1_G256_inv0;
    assign a1_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 = !axorb_1_G4_mul0_G16_mul1_G256_inv0;
    assign z5289_assgn5289 = r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    assign u0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (a0_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 & z1711_assgn1711);
    assign z5293_assgn5293 = r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    assign u1_hpc20_G4_mul0_G16_mul1_G256_inv0 = (a1_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 & z1713_assgn1713);
    assign v0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G4_mul0_G16_mul1_G256_inv0_reg ^ r0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign v1_hpc20_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G4_mul0_G16_mul1_G256_inv0_reg ^ r0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5301_assgn5301 = cxord_0_G4_mul0_G16_mul1_G256_inv0;
    assign p0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1719_assgn1719);
    assign p1_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & v1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p01_hpc20_G4_mul0_G16_mul1_G256_inv0 = (u0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul1_G256_inv0 = (p0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p01_hpc20_G4_mul0_G16_mul1_G256_inv0);
    assign z5311_assgn5311 = cxord_1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1727_assgn1727);
    assign p3_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & v0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p23_hpc20_G4_mul0_G16_mul1_G256_inv0 = (u1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p3_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p23_hpc20_G4_mul0_G16_mul1_G256_inv0);
    assign z5321_assgn5321 = dec_2_inp;
    assign r0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % z1735_assgn1735);
    assign a0_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 = !a0_G4_mul0_G16_mul1_G256_inv0;
    assign a1_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 = !a1_G4_mul0_G16_mul1_G256_inv0;
    assign z5329_assgn5329 = r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    assign u0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a0_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 & z1741_assgn1741);
    assign z5333_assgn5333 = r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    assign u1_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a1_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 & z1743_assgn1743);
    assign z5337_assgn5337 = c0_G4_mul0_G16_mul1_G256_inv0;
    assign v0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (z1746_assgn1746 ^ r0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5341_assgn5341 = c1_G4_mul0_G16_mul1_G256_inv0;
    assign v1_hpc21_G4_mul0_G16_mul1_G256_inv0 = (z1748_assgn1748 ^ r0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5345_assgn5345 = c0_G4_mul0_G16_mul1_G256_inv0;
    assign p0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1749_assgn1749);
    assign p1_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & v1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p01_hpc21_G4_mul0_G16_mul1_G256_inv0 = (u0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (p0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p01_hpc21_G4_mul0_G16_mul1_G256_inv0);
    assign z5355_assgn5355 = c1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1757_assgn1757);
    assign p3_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & v0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p23_hpc21_G4_mul0_G16_mul1_G256_inv0 = (u1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p3_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p23_hpc21_G4_mul0_G16_mul1_G256_inv0);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_G4_mul0_G16_mul1_G256_inv0 = (p1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign z5369_assgn5369 = dec_2_inp;
    assign r0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % z1769_assgn1769);
    assign a0_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 = !b0_G4_mul0_G16_mul1_G256_inv0;
    assign a1_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 = !b1_G4_mul0_G16_mul1_G256_inv0;
    assign z5377_assgn5377 = r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    assign u0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (a0_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 & z1775_assgn1775);
    assign z5381_assgn5381 = r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    assign u1_hpc22_G4_mul0_G16_mul1_G256_inv0 = (a1_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 & z1777_assgn1777);
    assign z5385_assgn5385 = d0_G4_mul0_G16_mul1_G256_inv0;
    assign v0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (z1780_assgn1780 ^ r0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5389_assgn5389 = d1_G4_mul0_G16_mul1_G256_inv0;
    assign v1_hpc22_G4_mul0_G16_mul1_G256_inv0 = (z1782_assgn1782 ^ r0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5393_assgn5393 = d0_G4_mul0_G16_mul1_G256_inv0;
    assign p0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1783_assgn1783);
    assign p1_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & v1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p01_hpc22_G4_mul0_G16_mul1_G256_inv0 = (u0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (p0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p01_hpc22_G4_mul0_G16_mul1_G256_inv0);
    assign z5403_assgn5403 = d1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1791_assgn1791);
    assign p3_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & v0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p23_hpc22_G4_mul0_G16_mul1_G256_inv0 = (u1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p3_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p23_hpc22_G4_mul0_G16_mul1_G256_inv0);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q1_G4_mul0_G16_mul1_G256_inv0 = (q1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign z5417_assgn5417 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul1_G256_inv0 = (p1_G4_mul0_G16_mul1_G256_inv0 << z1803_assgn1803);
    assign z5421_assgn5421 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << z1805_assgn1805);
    assign e0_G16_mul1_G256_inv0 = (p1ls1_G4_mul0_G16_mul1_G256_inv0 | q1_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign z5429_assgn5429 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1811_assgn1811);
    assign z5433_assgn5433 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1813_assgn1813);
    assign z5437_assgn5437 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1815_assgn1815);
    assign z5441_assgn5441 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1817_assgn1817);
    assign z5445_assgn5445 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1819_assgn1819);
    assign z5449_assgn5449 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1821_assgn1821);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign p1_G4_scl_N0_G16_mul1_G256_inv0 = b1_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign q1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_G4_scl_N0_G16_mul1_G256_inv0 ^ b1_G4_scl_N0_G16_mul1_G256_inv0);
    assign z5461_assgn5461 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p1_G4_scl_N0_G16_mul1_G256_inv0 << z1831_assgn1831);
    assign z5465_assgn5465 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << z1833_assgn1833);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign e11_G16_mul1_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul1_G256_inv0 | q1_G4_scl_N0_G16_mul1_G256_inv0);
    assign z5473_assgn5473 = z3_assgn3;
    assign r00_G4_mul1_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % z1839_assgn1839);
    assign z5477_assgn5477 = z3_assgn3;
    assign r10_G4_mul1_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % z1841_assgn1841);
    assign z5481_assgn5481 = z3_assgn3;
    assign r20_G4_mul1_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % z1843_assgn1843);
    assign z5485_assgn5485 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1845_assgn1845);
    assign z5489_assgn5489 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1847_assgn1847);
    assign z5493_assgn5493 = dec_1_inp;
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> z1849_assgn1849);
    assign z5497_assgn5497 = dec_1_inp;
    assign a1_G4_mul1_G16_mul1_G256_inv0 = (a1_0_G4_mul1_G16_mul1_G256_inv0 >> z1851_assgn1851);
    assign z5501_assgn5501 = dec_1_inp;
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1853_assgn1853);
    assign z5505_assgn5505 = dec_1_inp;
    assign b1_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1855_assgn1855);
    assign z5509_assgn5509 = dec_2_inp;
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & z1857_assgn1857);
    assign z5513_assgn5513 = dec_2_inp;
    assign c1_0_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & z1859_assgn1859);
    assign z5517_assgn5517 = dec_1_inp;
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> z1861_assgn1861);
    assign z5521_assgn5521 = dec_1_inp;
    assign c1_G4_mul1_G16_mul1_G256_inv0 = (c1_0_G4_mul1_G16_mul1_G256_inv0 >> z1863_assgn1863);
    assign z5525_assgn5525 = dec_1_inp;
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & z1865_assgn1865);
    assign z5529_assgn5529 = dec_1_inp;
    assign d1_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & z1867_assgn1867);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0_reg ^ d0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign axorb_1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ b1_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0_reg ^ d1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z5541_assgn5541 = dec_2_inp;
    assign r0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % z1877_assgn1877);
    assign a0_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 = !axorb_0_G4_mul1_G16_mul1_G256_inv0;
    assign a1_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 = !axorb_1_G4_mul1_G16_mul1_G256_inv0;
    assign z5549_assgn5549 = r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    assign u0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (a0_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 & z1883_assgn1883);
    assign z5553_assgn5553 = r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    assign u1_hpc20_G4_mul1_G16_mul1_G256_inv0 = (a1_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 & z1885_assgn1885);
    assign v0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (cxord_0_G4_mul1_G16_mul1_G256_inv0_reg ^ r0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign v1_hpc20_G4_mul1_G16_mul1_G256_inv0 = (cxord_1_G4_mul1_G16_mul1_G256_inv0_reg ^ r0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z5561_assgn5561 = cxord_0_G4_mul1_G16_mul1_G256_inv0;
    assign p0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1891_assgn1891);
    assign p1_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & v1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p01_hpc20_G4_mul1_G16_mul1_G256_inv0 = (u0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul1_G256_inv0 = (p0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p01_hpc20_G4_mul1_G16_mul1_G256_inv0);
    assign z5571_assgn5571 = cxord_1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1899_assgn1899);
    assign p3_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & v0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p23_hpc20_G4_mul1_G16_mul1_G256_inv0 = (u1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p3_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p23_hpc20_G4_mul1_G16_mul1_G256_inv0);
    assign z5581_assgn5581 = dec_2_inp;
    assign r0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % z1907_assgn1907);
    assign a0_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 = !a0_G4_mul1_G16_mul1_G256_inv0;
    assign a1_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 = !a1_G4_mul1_G16_mul1_G256_inv0;
    assign z5589_assgn5589 = r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    assign u0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a0_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 & z1913_assgn1913);
    assign z5593_assgn5593 = r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    assign u1_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a1_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 & z1915_assgn1915);
    assign z5597_assgn5597 = c0_G4_mul1_G16_mul1_G256_inv0;
    assign v0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (z1918_assgn1918 ^ r0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z5601_assgn5601 = c1_G4_mul1_G16_mul1_G256_inv0;
    assign v1_hpc21_G4_mul1_G16_mul1_G256_inv0 = (z1920_assgn1920 ^ r0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z5605_assgn5605 = c0_G4_mul1_G16_mul1_G256_inv0;
    assign p0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1921_assgn1921);
    assign p1_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & v1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p01_hpc21_G4_mul1_G16_mul1_G256_inv0 = (u0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (p0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p01_hpc21_G4_mul1_G16_mul1_G256_inv0);
    assign z5615_assgn5615 = c1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1929_assgn1929);
    assign p3_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & v0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p23_hpc21_G4_mul1_G16_mul1_G256_inv0 = (u1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p3_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p23_hpc21_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_G4_mul1_G16_mul1_G256_inv0 = (p1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign z5629_assgn5629 = dec_2_inp;
    assign r0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % z1941_assgn1941);
    assign a0_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 = !b0_G4_mul1_G16_mul1_G256_inv0;
    assign a1_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 = !b1_G4_mul1_G16_mul1_G256_inv0;
    assign z5637_assgn5637 = r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    assign u0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (a0_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 & z1947_assgn1947);
    assign z5641_assgn5641 = r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    assign u1_hpc22_G4_mul1_G16_mul1_G256_inv0 = (a1_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 & z1949_assgn1949);
    assign z5645_assgn5645 = d0_G4_mul1_G16_mul1_G256_inv0;
    assign v0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (z1952_assgn1952 ^ r0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z5649_assgn5649 = d1_G4_mul1_G16_mul1_G256_inv0;
    assign v1_hpc22_G4_mul1_G16_mul1_G256_inv0 = (z1954_assgn1954 ^ r0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z5653_assgn5653 = d0_G4_mul1_G16_mul1_G256_inv0;
    assign p0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1955_assgn1955);
    assign p1_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & v1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p01_hpc22_G4_mul1_G16_mul1_G256_inv0 = (u0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (p0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p01_hpc22_G4_mul1_G16_mul1_G256_inv0);
    assign z5663_assgn5663 = d1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1963_assgn1963);
    assign p3_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & v0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p23_hpc22_G4_mul1_G16_mul1_G256_inv0 = (u1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p3_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p23_hpc22_G4_mul1_G16_mul1_G256_inv0);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q1_G4_mul1_G16_mul1_G256_inv0 = (q1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign z5677_assgn5677 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul1_G256_inv0 = (p1_G4_mul1_G16_mul1_G256_inv0 << z1975_assgn1975);
    assign z5681_assgn5681 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << z1977_assgn1977);
    assign p0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul1_G16_mul1_G256_inv0 | q1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p1_G16_mul1_G256_inv0 = (p1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign z5693_assgn5693 = z3_assgn3;
    assign r00_G4_mul2_G16_mul1_G256_inv0 = (r60_G16_mul1_G256_inv0 % z1987_assgn1987);
    assign z5697_assgn5697 = z3_assgn3;
    assign r10_G4_mul2_G16_mul1_G256_inv0 = (r70_G16_mul1_G256_inv0 % z1989_assgn1989);
    assign z5701_assgn5701 = z3_assgn3;
    assign r20_G4_mul2_G16_mul1_G256_inv0 = (r80_G16_mul1_G256_inv0 % z1991_assgn1991);
    assign z5705_assgn5705 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1993_assgn1993);
    assign z5709_assgn5709 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1995_assgn1995);
    assign z5713_assgn5713 = dec_1_inp;
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> z1997_assgn1997);
    assign z5717_assgn5717 = dec_1_inp;
    assign a1_G4_mul2_G16_mul1_G256_inv0 = (a1_0_G4_mul2_G16_mul1_G256_inv0 >> z1999_assgn1999);
    assign z5721_assgn5721 = dec_1_inp;
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z2001_assgn2001);
    assign z5725_assgn5725 = dec_1_inp;
    assign b1_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z2003_assgn2003);
    assign z5729_assgn5729 = dec_2_inp;
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & z2005_assgn2005);
    assign z5733_assgn5733 = dec_2_inp;
    assign c1_0_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & z2007_assgn2007);
    assign z5737_assgn5737 = dec_1_inp;
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> z2009_assgn2009);
    assign z5741_assgn5741 = dec_1_inp;
    assign c1_G4_mul2_G16_mul1_G256_inv0 = (c1_0_G4_mul2_G16_mul1_G256_inv0 >> z2011_assgn2011);
    assign z5745_assgn5745 = dec_1_inp;
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & z2013_assgn2013);
    assign z5749_assgn5749 = dec_1_inp;
    assign d1_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & z2015_assgn2015);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0_reg ^ d0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign axorb_1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ b1_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0_reg ^ d1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z5761_assgn5761 = dec_2_inp;
    assign r0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % z2025_assgn2025);
    assign a0_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 = !axorb_0_G4_mul2_G16_mul1_G256_inv0;
    assign a1_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 = !axorb_1_G4_mul2_G16_mul1_G256_inv0;
    assign z5769_assgn5769 = r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    assign u0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (a0_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 & z2031_assgn2031);
    assign z5773_assgn5773 = r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    assign u1_hpc20_G4_mul2_G16_mul1_G256_inv0 = (a1_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 & z2033_assgn2033);
    assign v0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (cxord_0_G4_mul2_G16_mul1_G256_inv0_reg ^ r0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign v1_hpc20_G4_mul2_G16_mul1_G256_inv0 = (cxord_1_G4_mul2_G16_mul1_G256_inv0_reg ^ r0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z5781_assgn5781 = cxord_0_G4_mul2_G16_mul1_G256_inv0;
    assign p0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z2039_assgn2039);
    assign p1_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & v1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p01_hpc20_G4_mul2_G16_mul1_G256_inv0 = (u0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul1_G256_inv0 = (p0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p01_hpc20_G4_mul2_G16_mul1_G256_inv0);
    assign z5791_assgn5791 = cxord_1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z2047_assgn2047);
    assign p3_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & v0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p23_hpc20_G4_mul2_G16_mul1_G256_inv0 = (u1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p3_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p23_hpc20_G4_mul2_G16_mul1_G256_inv0);
    assign z5801_assgn5801 = dec_2_inp;
    assign r0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % z2055_assgn2055);
    assign a0_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 = !a0_G4_mul2_G16_mul1_G256_inv0;
    assign a1_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 = !a1_G4_mul2_G16_mul1_G256_inv0;
    assign z5809_assgn5809 = r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    assign u0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a0_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 & z2061_assgn2061);
    assign z5813_assgn5813 = r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    assign u1_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a1_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 & z2063_assgn2063);
    assign z5817_assgn5817 = c0_G4_mul2_G16_mul1_G256_inv0;
    assign v0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (z2066_assgn2066 ^ r0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z5821_assgn5821 = c1_G4_mul2_G16_mul1_G256_inv0;
    assign v1_hpc21_G4_mul2_G16_mul1_G256_inv0 = (z2068_assgn2068 ^ r0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z5825_assgn5825 = c0_G4_mul2_G16_mul1_G256_inv0;
    assign p0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z2069_assgn2069);
    assign p1_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & v1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p01_hpc21_G4_mul2_G16_mul1_G256_inv0 = (u0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (p0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p01_hpc21_G4_mul2_G16_mul1_G256_inv0);
    assign z5835_assgn5835 = c1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z2077_assgn2077);
    assign p3_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & v0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p23_hpc21_G4_mul2_G16_mul1_G256_inv0 = (u1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p3_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p23_hpc21_G4_mul2_G16_mul1_G256_inv0);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_G4_mul2_G16_mul1_G256_inv0 = (p1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign z5849_assgn5849 = dec_2_inp;
    assign r0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % z2089_assgn2089);
    assign a0_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 = !b0_G4_mul2_G16_mul1_G256_inv0;
    assign a1_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 = !b1_G4_mul2_G16_mul1_G256_inv0;
    assign z5857_assgn5857 = r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    assign u0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (a0_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 & z2095_assgn2095);
    assign z5861_assgn5861 = r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    assign u1_hpc22_G4_mul2_G16_mul1_G256_inv0 = (a1_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 & z2097_assgn2097);
    assign z5865_assgn5865 = d0_G4_mul2_G16_mul1_G256_inv0;
    assign v0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (z2100_assgn2100 ^ r0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z5869_assgn5869 = d1_G4_mul2_G16_mul1_G256_inv0;
    assign v1_hpc22_G4_mul2_G16_mul1_G256_inv0 = (z2102_assgn2102 ^ r0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z5873_assgn5873 = d0_G4_mul2_G16_mul1_G256_inv0;
    assign p0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z2103_assgn2103);
    assign p1_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & v1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p01_hpc22_G4_mul2_G16_mul1_G256_inv0 = (u0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (p0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p01_hpc22_G4_mul2_G16_mul1_G256_inv0);
    assign z5883_assgn5883 = d1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z2111_assgn2111);
    assign p3_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & v0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p23_hpc22_G4_mul2_G16_mul1_G256_inv0 = (u1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p3_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p23_hpc22_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q1_G4_mul2_G16_mul1_G256_inv0 = (q1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign z5897_assgn5897 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul1_G256_inv0 = (p1_G4_mul2_G16_mul1_G256_inv0 << z2123_assgn2123);
    assign z5901_assgn5901 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << z2125_assgn2125);
    assign q0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul2_G16_mul1_G256_inv0 | q1_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign q1_G16_mul1_G256_inv0 = (q1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign z5913_assgn5913 = dec_2_inp;
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << z2135_assgn2135);
    assign z5917_assgn5917 = dec_2_inp;
    assign p1ls2_G16_mul1_G256_inv0 = (p1_G16_mul1_G256_inv0 << z2137_assgn2137);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign p1_G256_inv0 = (p1ls2_G16_mul1_G256_inv0 | q1_G16_mul1_G256_inv0);
    assign z5925_assgn5925 = z1_assgn1;
    assign r00_G16_mul2_G256_inv0 = (r27_inp % z2143_assgn2143);
    assign z5929_assgn5929 = z1_assgn1;
    assign r10_G16_mul2_G256_inv0 = (r28_inp % z2145_assgn2145);
    assign z5933_assgn5933 = z1_assgn1;
    assign r20_G16_mul2_G256_inv0 = (r29_inp % z2147_assgn2147);
    assign z5937_assgn5937 = z1_assgn1;
    assign r30_G16_mul2_G256_inv0 = (r30_inp % z2149_assgn2149);
    assign z5941_assgn5941 = z1_assgn1;
    assign r40_G16_mul2_G256_inv0 = (r31_inp % z2151_assgn2151);
    assign z5945_assgn5945 = z1_assgn1;
    assign r50_G16_mul2_G256_inv0 = (r32_inp % z2153_assgn2153);
    assign z5949_assgn5949 = z1_assgn1;
    assign r60_G16_mul2_G256_inv0 = (r33_inp % z2155_assgn2155);
    assign z5953_assgn5953 = z1_assgn1;
    assign r70_G16_mul2_G256_inv0 = (r34_inp % z2157_assgn2157);
    assign z5957_assgn5957 = z1_assgn1;
    assign r80_G16_mul2_G256_inv0 = (r35_inp % z2159_assgn2159);
    assign z5961_assgn5961 = dec_12_inp;
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z2161_assgn2161);
    assign z5965_assgn5965 = dec_12_inp;
    assign a1_0_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2163_assgn2163);
    assign z5969_assgn5969 = dec_2_inp;
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> z2165_assgn2165);
    assign z5973_assgn5973 = dec_2_inp;
    assign a1_G16_mul2_G256_inv0 = (a1_0_G16_mul2_G256_inv0 >> z2167_assgn2167);
    assign z5977_assgn5977 = dec_3_inp;
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z2169_assgn2169);
    assign z5981_assgn5981 = dec_3_inp;
    assign b1_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2171_assgn2171);
    assign z5985_assgn5985 = dec_12_inp;
    assign z5987_assgn5987 = a0_G256_inv0;
    assign c0_0_G16_mul2_G256_inv0 = (z2174_assgn2174 & z2173_assgn2173);
    assign z5991_assgn5991 = dec_12_inp;
    assign z5993_assgn5993 = a1_G256_inv0;
    assign c1_0_G16_mul2_G256_inv0 = (z2176_assgn2176 & z2175_assgn2175);
    assign z5997_assgn5997 = dec_2_inp;
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> z2177_assgn2177);
    assign z6001_assgn6001 = dec_2_inp;
    assign c1_G16_mul2_G256_inv0 = (c1_0_G16_mul2_G256_inv0 >> z2179_assgn2179);
    assign z6005_assgn6005 = dec_3_inp;
    assign z6007_assgn6007 = a0_G256_inv0;
    assign d0_G16_mul2_G256_inv0 = (z2182_assgn2182 & z2181_assgn2181);
    assign z6011_assgn6011 = dec_3_inp;
    assign z6013_assgn6013 = a1_G256_inv0;
    assign d1_G16_mul2_G256_inv0 = (z2184_assgn2184 & z2183_assgn2183);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign axorb_1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 ^ b1_G16_mul2_G256_inv0);
    assign cxord_1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 ^ d1_G16_mul2_G256_inv0);
    assign z6025_assgn6025 = z3_assgn3;
    assign r00_G4_mul0_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % z2193_assgn2193);
    assign z6029_assgn6029 = z3_assgn3;
    assign r10_G4_mul0_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % z2195_assgn2195);
    assign z6033_assgn6033 = z3_assgn3;
    assign r20_G4_mul0_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % z2197_assgn2197);
    assign z6037_assgn6037 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z2199_assgn2199);
    assign z6041_assgn6041 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2201_assgn2201);
    assign z6045_assgn6045 = dec_1_inp;
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> z2203_assgn2203);
    assign z6049_assgn6049 = dec_1_inp;
    assign a1_G4_mul0_G16_mul2_G256_inv0 = (a1_0_G4_mul0_G16_mul2_G256_inv0 >> z2205_assgn2205);
    assign z6053_assgn6053 = dec_1_inp;
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z2207_assgn2207);
    assign z6057_assgn6057 = dec_1_inp;
    assign b1_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2209_assgn2209);
    assign z6061_assgn6061 = dec_2_inp;
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & z2211_assgn2211);
    assign z6065_assgn6065 = dec_2_inp;
    assign c1_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & z2213_assgn2213);
    assign z6069_assgn6069 = dec_1_inp;
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> z2215_assgn2215);
    assign z6073_assgn6073 = dec_1_inp;
    assign c1_G4_mul0_G16_mul2_G256_inv0 = (c1_0_G4_mul0_G16_mul2_G256_inv0 >> z2217_assgn2217);
    assign z6077_assgn6077 = dec_1_inp;
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & z2219_assgn2219);
    assign z6081_assgn6081 = dec_1_inp;
    assign d1_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & z2221_assgn2221);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0_reg ^ d0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign axorb_1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ b1_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0_reg ^ d1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6093_assgn6093 = dec_2_inp;
    assign r0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % z2231_assgn2231);
    assign a0_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 = !axorb_0_G4_mul0_G16_mul2_G256_inv0;
    assign a1_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 = !axorb_1_G4_mul0_G16_mul2_G256_inv0;
    assign z6101_assgn6101 = r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    assign u0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (a0_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 & z2237_assgn2237);
    assign z6105_assgn6105 = r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    assign u1_hpc20_G4_mul0_G16_mul2_G256_inv0 = (a1_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 & z2239_assgn2239);
    assign v0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G4_mul0_G16_mul2_G256_inv0_reg ^ r0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign v1_hpc20_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G4_mul0_G16_mul2_G256_inv0_reg ^ r0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6113_assgn6113 = cxord_0_G4_mul0_G16_mul2_G256_inv0;
    assign p0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z2245_assgn2245);
    assign p1_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & v1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p01_hpc20_G4_mul0_G16_mul2_G256_inv0 = (u0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul2_G256_inv0 = (p0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p01_hpc20_G4_mul0_G16_mul2_G256_inv0);
    assign z6123_assgn6123 = cxord_1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z2253_assgn2253);
    assign p3_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & v0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p23_hpc20_G4_mul0_G16_mul2_G256_inv0 = (u1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p3_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p23_hpc20_G4_mul0_G16_mul2_G256_inv0);
    assign z6133_assgn6133 = dec_2_inp;
    assign r0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % z2261_assgn2261);
    assign a0_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 = !a0_G4_mul0_G16_mul2_G256_inv0;
    assign a1_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 = !a1_G4_mul0_G16_mul2_G256_inv0;
    assign z6141_assgn6141 = r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    assign u0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a0_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 & z2267_assgn2267);
    assign z6145_assgn6145 = r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    assign u1_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a1_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 & z2269_assgn2269);
    assign z6149_assgn6149 = c0_G4_mul0_G16_mul2_G256_inv0;
    assign v0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (z2272_assgn2272 ^ r0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6153_assgn6153 = c1_G4_mul0_G16_mul2_G256_inv0;
    assign v1_hpc21_G4_mul0_G16_mul2_G256_inv0 = (z2274_assgn2274 ^ r0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6157_assgn6157 = c0_G4_mul0_G16_mul2_G256_inv0;
    assign p0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z2275_assgn2275);
    assign p1_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & v1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p01_hpc21_G4_mul0_G16_mul2_G256_inv0 = (u0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul2_G256_inv0 = (p0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p01_hpc21_G4_mul0_G16_mul2_G256_inv0);
    assign z6167_assgn6167 = c1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z2283_assgn2283);
    assign p3_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & v0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p23_hpc21_G4_mul0_G16_mul2_G256_inv0 = (u1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p3_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p23_hpc21_G4_mul0_G16_mul2_G256_inv0);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_G4_mul0_G16_mul2_G256_inv0 = (p1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign z6181_assgn6181 = dec_2_inp;
    assign r0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % z2295_assgn2295);
    assign a0_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 = !b0_G4_mul0_G16_mul2_G256_inv0;
    assign a1_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 = !b1_G4_mul0_G16_mul2_G256_inv0;
    assign z6189_assgn6189 = r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    assign u0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (a0_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 & z2301_assgn2301);
    assign z6193_assgn6193 = r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    assign u1_hpc22_G4_mul0_G16_mul2_G256_inv0 = (a1_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 & z2303_assgn2303);
    assign z6197_assgn6197 = d0_G4_mul0_G16_mul2_G256_inv0;
    assign v0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (z2306_assgn2306 ^ r0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6201_assgn6201 = d1_G4_mul0_G16_mul2_G256_inv0;
    assign v1_hpc22_G4_mul0_G16_mul2_G256_inv0 = (z2308_assgn2308 ^ r0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6205_assgn6205 = d0_G4_mul0_G16_mul2_G256_inv0;
    assign p0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z2309_assgn2309);
    assign p1_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & v1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p01_hpc22_G4_mul0_G16_mul2_G256_inv0 = (u0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul2_G256_inv0 = (p0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p01_hpc22_G4_mul0_G16_mul2_G256_inv0);
    assign z6215_assgn6215 = d1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z2317_assgn2317);
    assign p3_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & v0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p23_hpc22_G4_mul0_G16_mul2_G256_inv0 = (u1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p3_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p23_hpc22_G4_mul0_G16_mul2_G256_inv0);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q1_G4_mul0_G16_mul2_G256_inv0 = (q1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign z6229_assgn6229 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul2_G256_inv0 = (p1_G4_mul0_G16_mul2_G256_inv0 << z2329_assgn2329);
    assign z6233_assgn6233 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << z2331_assgn2331);
    assign e0_G16_mul2_G256_inv0 = (p1ls1_G4_mul0_G16_mul2_G256_inv0 | q1_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign z6241_assgn6241 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z2337_assgn2337);
    assign z6245_assgn6245 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2339_assgn2339);
    assign z6249_assgn6249 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2341_assgn2341);
    assign z6253_assgn6253 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2343_assgn2343);
    assign z6257_assgn6257 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z2345_assgn2345);
    assign z6261_assgn6261 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2347_assgn2347);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign p1_G4_scl_N0_G16_mul2_G256_inv0 = b1_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign q1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_G4_scl_N0_G16_mul2_G256_inv0 ^ b1_G4_scl_N0_G16_mul2_G256_inv0);
    assign z6273_assgn6273 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p1_G4_scl_N0_G16_mul2_G256_inv0 << z2357_assgn2357);
    assign z6277_assgn6277 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << z2359_assgn2359);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign e11_G16_mul2_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul2_G256_inv0 | q1_G4_scl_N0_G16_mul2_G256_inv0);
    assign z6285_assgn6285 = z3_assgn3;
    assign r00_G4_mul1_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % z2365_assgn2365);
    assign z6289_assgn6289 = z3_assgn3;
    assign r10_G4_mul1_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % z2367_assgn2367);
    assign z6293_assgn6293 = z3_assgn3;
    assign r20_G4_mul1_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % z2369_assgn2369);
    assign z6297_assgn6297 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z2371_assgn2371);
    assign z6301_assgn6301 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2373_assgn2373);
    assign z6305_assgn6305 = dec_1_inp;
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> z2375_assgn2375);
    assign z6309_assgn6309 = dec_1_inp;
    assign a1_G4_mul1_G16_mul2_G256_inv0 = (a1_0_G4_mul1_G16_mul2_G256_inv0 >> z2377_assgn2377);
    assign z6313_assgn6313 = dec_1_inp;
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z2379_assgn2379);
    assign z6317_assgn6317 = dec_1_inp;
    assign b1_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2381_assgn2381);
    assign z6321_assgn6321 = dec_2_inp;
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & z2383_assgn2383);
    assign z6325_assgn6325 = dec_2_inp;
    assign c1_0_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & z2385_assgn2385);
    assign z6329_assgn6329 = dec_1_inp;
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> z2387_assgn2387);
    assign z6333_assgn6333 = dec_1_inp;
    assign c1_G4_mul1_G16_mul2_G256_inv0 = (c1_0_G4_mul1_G16_mul2_G256_inv0 >> z2389_assgn2389);
    assign z6337_assgn6337 = dec_1_inp;
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & z2391_assgn2391);
    assign z6341_assgn6341 = dec_1_inp;
    assign d1_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & z2393_assgn2393);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0_reg ^ d0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign axorb_1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ b1_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0_reg ^ d1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z6353_assgn6353 = dec_2_inp;
    assign r0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % z2403_assgn2403);
    assign a0_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 = !axorb_0_G4_mul1_G16_mul2_G256_inv0;
    assign a1_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 = !axorb_1_G4_mul1_G16_mul2_G256_inv0;
    assign z6361_assgn6361 = r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    assign u0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (a0_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 & z2409_assgn2409);
    assign z6365_assgn6365 = r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    assign u1_hpc20_G4_mul1_G16_mul2_G256_inv0 = (a1_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 & z2411_assgn2411);
    assign v0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (cxord_0_G4_mul1_G16_mul2_G256_inv0_reg ^ r0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign v1_hpc20_G4_mul1_G16_mul2_G256_inv0 = (cxord_1_G4_mul1_G16_mul2_G256_inv0_reg ^ r0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z6373_assgn6373 = cxord_0_G4_mul1_G16_mul2_G256_inv0;
    assign p0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2417_assgn2417);
    assign p1_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & v1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p01_hpc20_G4_mul1_G16_mul2_G256_inv0 = (u0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul2_G256_inv0 = (p0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p01_hpc20_G4_mul1_G16_mul2_G256_inv0);
    assign z6383_assgn6383 = cxord_1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2425_assgn2425);
    assign p3_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & v0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p23_hpc20_G4_mul1_G16_mul2_G256_inv0 = (u1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p3_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p23_hpc20_G4_mul1_G16_mul2_G256_inv0);
    assign z6393_assgn6393 = dec_2_inp;
    assign r0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % z2433_assgn2433);
    assign a0_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 = !a0_G4_mul1_G16_mul2_G256_inv0;
    assign a1_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 = !a1_G4_mul1_G16_mul2_G256_inv0;
    assign z6401_assgn6401 = r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    assign u0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a0_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 & z2439_assgn2439);
    assign z6405_assgn6405 = r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    assign u1_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a1_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 & z2441_assgn2441);
    assign z6409_assgn6409 = c0_G4_mul1_G16_mul2_G256_inv0;
    assign v0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (z2444_assgn2444 ^ r0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z6413_assgn6413 = c1_G4_mul1_G16_mul2_G256_inv0;
    assign v1_hpc21_G4_mul1_G16_mul2_G256_inv0 = (z2446_assgn2446 ^ r0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z6417_assgn6417 = c0_G4_mul1_G16_mul2_G256_inv0;
    assign p0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2447_assgn2447);
    assign p1_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & v1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p01_hpc21_G4_mul1_G16_mul2_G256_inv0 = (u0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul2_G256_inv0 = (p0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p01_hpc21_G4_mul1_G16_mul2_G256_inv0);
    assign z6427_assgn6427 = c1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2455_assgn2455);
    assign p3_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & v0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p23_hpc21_G4_mul1_G16_mul2_G256_inv0 = (u1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p3_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p23_hpc21_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_G4_mul1_G16_mul2_G256_inv0 = (p1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign z6441_assgn6441 = dec_2_inp;
    assign r0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % z2467_assgn2467);
    assign a0_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 = !b0_G4_mul1_G16_mul2_G256_inv0;
    assign a1_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 = !b1_G4_mul1_G16_mul2_G256_inv0;
    assign z6449_assgn6449 = r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    assign u0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (a0_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 & z2473_assgn2473);
    assign z6453_assgn6453 = r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    assign u1_hpc22_G4_mul1_G16_mul2_G256_inv0 = (a1_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 & z2475_assgn2475);
    assign z6457_assgn6457 = d0_G4_mul1_G16_mul2_G256_inv0;
    assign v0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (z2478_assgn2478 ^ r0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z6461_assgn6461 = d1_G4_mul1_G16_mul2_G256_inv0;
    assign v1_hpc22_G4_mul1_G16_mul2_G256_inv0 = (z2480_assgn2480 ^ r0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z6465_assgn6465 = d0_G4_mul1_G16_mul2_G256_inv0;
    assign p0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2481_assgn2481);
    assign p1_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & v1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p01_hpc22_G4_mul1_G16_mul2_G256_inv0 = (u0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul2_G256_inv0 = (p0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p01_hpc22_G4_mul1_G16_mul2_G256_inv0);
    assign z6475_assgn6475 = d1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2489_assgn2489);
    assign p3_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & v0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p23_hpc22_G4_mul1_G16_mul2_G256_inv0 = (u1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p3_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p23_hpc22_G4_mul1_G16_mul2_G256_inv0);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q1_G4_mul1_G16_mul2_G256_inv0 = (q1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign z6489_assgn6489 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul2_G256_inv0 = (p1_G4_mul1_G16_mul2_G256_inv0 << z2501_assgn2501);
    assign z6493_assgn6493 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << z2503_assgn2503);
    assign p0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul1_G16_mul2_G256_inv0 | q1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p1_G16_mul2_G256_inv0 = (p1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign z6505_assgn6505 = z3_assgn3;
    assign r00_G4_mul2_G16_mul2_G256_inv0 = (r60_G16_mul2_G256_inv0 % z2513_assgn2513);
    assign z6509_assgn6509 = z3_assgn3;
    assign r10_G4_mul2_G16_mul2_G256_inv0 = (r70_G16_mul2_G256_inv0 % z2515_assgn2515);
    assign z6513_assgn6513 = z3_assgn3;
    assign r20_G4_mul2_G16_mul2_G256_inv0 = (r80_G16_mul2_G256_inv0 % z2517_assgn2517);
    assign z6517_assgn6517 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2519_assgn2519);
    assign z6521_assgn6521 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2521_assgn2521);
    assign z6525_assgn6525 = dec_1_inp;
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> z2523_assgn2523);
    assign z6529_assgn6529 = dec_1_inp;
    assign a1_G4_mul2_G16_mul2_G256_inv0 = (a1_0_G4_mul2_G16_mul2_G256_inv0 >> z2525_assgn2525);
    assign z6533_assgn6533 = dec_1_inp;
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2527_assgn2527);
    assign z6537_assgn6537 = dec_1_inp;
    assign b1_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2529_assgn2529);
    assign z6541_assgn6541 = dec_2_inp;
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & z2531_assgn2531);
    assign z6545_assgn6545 = dec_2_inp;
    assign c1_0_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & z2533_assgn2533);
    assign z6549_assgn6549 = dec_1_inp;
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> z2535_assgn2535);
    assign z6553_assgn6553 = dec_1_inp;
    assign c1_G4_mul2_G16_mul2_G256_inv0 = (c1_0_G4_mul2_G16_mul2_G256_inv0 >> z2537_assgn2537);
    assign z6557_assgn6557 = dec_1_inp;
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & z2539_assgn2539);
    assign z6561_assgn6561 = dec_1_inp;
    assign d1_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & z2541_assgn2541);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0_reg ^ d0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign axorb_1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ b1_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0_reg ^ d1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z6573_assgn6573 = dec_2_inp;
    assign r0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % z2551_assgn2551);
    assign a0_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 = !axorb_0_G4_mul2_G16_mul2_G256_inv0;
    assign a1_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 = !axorb_1_G4_mul2_G16_mul2_G256_inv0;
    assign z6581_assgn6581 = r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    assign u0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (a0_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 & z2557_assgn2557);
    assign z6585_assgn6585 = r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    assign u1_hpc20_G4_mul2_G16_mul2_G256_inv0 = (a1_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 & z2559_assgn2559);
    assign v0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (cxord_0_G4_mul2_G16_mul2_G256_inv0_reg ^ r0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign v1_hpc20_G4_mul2_G16_mul2_G256_inv0 = (cxord_1_G4_mul2_G16_mul2_G256_inv0_reg ^ r0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z6593_assgn6593 = cxord_0_G4_mul2_G16_mul2_G256_inv0;
    assign p0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2565_assgn2565);
    assign p1_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & v1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p01_hpc20_G4_mul2_G16_mul2_G256_inv0 = (u0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul2_G256_inv0 = (p0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p01_hpc20_G4_mul2_G16_mul2_G256_inv0);
    assign z6603_assgn6603 = cxord_1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2573_assgn2573);
    assign p3_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & v0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p23_hpc20_G4_mul2_G16_mul2_G256_inv0 = (u1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p3_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p23_hpc20_G4_mul2_G16_mul2_G256_inv0);
    assign z6613_assgn6613 = dec_2_inp;
    assign r0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % z2581_assgn2581);
    assign a0_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 = !a0_G4_mul2_G16_mul2_G256_inv0;
    assign a1_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 = !a1_G4_mul2_G16_mul2_G256_inv0;
    assign z6621_assgn6621 = r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    assign u0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a0_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 & z2587_assgn2587);
    assign z6625_assgn6625 = r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    assign u1_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a1_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 & z2589_assgn2589);
    assign z6629_assgn6629 = c0_G4_mul2_G16_mul2_G256_inv0;
    assign v0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (z2592_assgn2592 ^ r0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z6633_assgn6633 = c1_G4_mul2_G16_mul2_G256_inv0;
    assign v1_hpc21_G4_mul2_G16_mul2_G256_inv0 = (z2594_assgn2594 ^ r0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z6637_assgn6637 = c0_G4_mul2_G16_mul2_G256_inv0;
    assign p0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2595_assgn2595);
    assign p1_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & v1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p01_hpc21_G4_mul2_G16_mul2_G256_inv0 = (u0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul2_G256_inv0 = (p0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p01_hpc21_G4_mul2_G16_mul2_G256_inv0);
    assign z6647_assgn6647 = c1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2603_assgn2603);
    assign p3_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & v0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p23_hpc21_G4_mul2_G16_mul2_G256_inv0 = (u1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p3_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p23_hpc21_G4_mul2_G16_mul2_G256_inv0);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_G4_mul2_G16_mul2_G256_inv0 = (p1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign z6661_assgn6661 = dec_2_inp;
    assign r0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % z2615_assgn2615);
    assign a0_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 = !b0_G4_mul2_G16_mul2_G256_inv0;
    assign a1_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 = !b1_G4_mul2_G16_mul2_G256_inv0;
    assign z6669_assgn6669 = r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    assign u0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (a0_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 & z2621_assgn2621);
    assign z6673_assgn6673 = r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    assign u1_hpc22_G4_mul2_G16_mul2_G256_inv0 = (a1_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 & z2623_assgn2623);
    assign z6677_assgn6677 = d0_G4_mul2_G16_mul2_G256_inv0;
    assign v0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (z2626_assgn2626 ^ r0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z6681_assgn6681 = d1_G4_mul2_G16_mul2_G256_inv0;
    assign v1_hpc22_G4_mul2_G16_mul2_G256_inv0 = (z2628_assgn2628 ^ r0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z6685_assgn6685 = d0_G4_mul2_G16_mul2_G256_inv0;
    assign p0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2629_assgn2629);
    assign p1_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & v1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p01_hpc22_G4_mul2_G16_mul2_G256_inv0 = (u0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul2_G256_inv0 = (p0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p01_hpc22_G4_mul2_G16_mul2_G256_inv0);
    assign z6695_assgn6695 = d1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2637_assgn2637);
    assign p3_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & v0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p23_hpc22_G4_mul2_G16_mul2_G256_inv0 = (u1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p3_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p23_hpc22_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q1_G4_mul2_G16_mul2_G256_inv0 = (q1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign z6709_assgn6709 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul2_G256_inv0 = (p1_G4_mul2_G16_mul2_G256_inv0 << z2649_assgn2649);
    assign z6713_assgn6713 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << z2651_assgn2651);
    assign q0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul2_G16_mul2_G256_inv0 | q1_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign q1_G16_mul2_G256_inv0 = (q1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign z6725_assgn6725 = dec_2_inp;
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << z2661_assgn2661);
    assign z6729_assgn6729 = dec_2_inp;
    assign p1ls2_G16_mul2_G256_inv0 = (p1_G16_mul2_G256_inv0 << z2663_assgn2663);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign q1_G256_inv0 = (p1ls2_G16_mul2_G256_inv0 | q1_G16_mul2_G256_inv0);
    assign z6737_assgn6737 = z3_assgn3;
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << z2669_assgn2669);
    assign z6741_assgn6741 = z3_assgn3;
    assign p1ls4_G256_inv0 = (p1_G256_inv0 << z2671_assgn2671);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign t5 = (p1ls4_G256_inv0 | q1_G256_inv0);
    assign z6749_assgn6749 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign z6753_assgn6753 = dec_1_inp;
    assign cond1_G256_newbasis1 = (t4 & z2681_assgn2681);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * yxorb1_G256_newbasis1);
    assign tempyIntoNegCond1_G256_newbasis1 = (tempy1_G256_newbasis1 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempyIntoNegCond1_G256_newbasis1);
    assign z6767_assgn6767 = dec_1_inp;
    assign x1_G256_newbasis1 = (t4 >> z2693_assgn2693);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign z6773_assgn6773 = dec_1_inp;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & z2697_assgn2697);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign z6779_assgn6779 = dec_3_inp;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ z2701_assgn2701);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempyIntoNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempyIntoNegCond2_G256_newbasis1);
    assign z6789_assgn6789 = dec_1_inp;
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> z2709_assgn2709);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign z6795_assgn6795 = dec_1_inp;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & z2713_assgn2713);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign z6801_assgn6801 = z3_assgn3;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ z2717_assgn2717);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempyIntoNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempyIntoNegCond3_G256_newbasis1);
    assign z6811_assgn6811 = dec_1_inp;
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> z2725_assgn2725);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign z6817_assgn6817 = dec_1_inp;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & z2729_assgn2729);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ dec_220_inp);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempyIntoNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempyIntoNegCond4_G256_newbasis1);
    assign z6831_assgn6831 = dec_1_inp;
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> z2741_assgn2741);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign z6837_assgn6837 = dec_1_inp;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & z2745_assgn2745);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ dec_11_inp);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempyIntoNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempyIntoNegCond5_G256_newbasis1);
    assign z6851_assgn6851 = dec_1_inp;
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> z2757_assgn2757);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign z6857_assgn6857 = dec_1_inp;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & z2761_assgn2761);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ dec_158_inp);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempyIntoNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempyIntoNegCond6_G256_newbasis1);
    assign z6871_assgn6871 = dec_1_inp;
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> z2773_assgn2773);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign z6877_assgn6877 = dec_1_inp;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & z2777_assgn2777);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ dec_45_inp);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempyIntoNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempyIntoNegCond7_G256_newbasis1);
    assign z6891_assgn6891 = dec_1_inp;
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> z2789_assgn2789);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign z6897_assgn6897 = dec_1_inp;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & z2793_assgn2793);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ dec_88_inp);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempyIntoNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempyIntoNegCond8_G256_newbasis1);
    assign z6911_assgn6911 = dec_1_inp;
    assign x8_G256_newbasis1 = (x7_G256_newbasis1 >> z2805_assgn2805);
    assign t6 = y8_G256_newbasis1;
    assign z6917_assgn6917 = dec_0_inp;
    assign z_tempy1_G256_newbasis1 = z_y_G256_newbasis1;
    assign z6921_assgn6921 = dec_1_inp;
    assign z_cond1_G256_newbasis1 = (t5 & z2813_assgn2813);
    assign z_negCond1_G256_newbasis1 = !z_cond1_G256_newbasis1;
    assign z_yxorb1_G256_newbasis1 = (z_y_G256_newbasis1 ^ dec_36_inp);
    assign z_ny1_G256_newbasis1 = (z_cond1_G256_newbasis1 * z_yxorb1_G256_newbasis1);
    assign z_tempyIntoNegCond1_G256_newbasis1 = (z_tempy1_G256_newbasis1 * z_negCond1_G256_newbasis1);
    assign z_y1_G256_newbasis1 = (z_ny1_G256_newbasis1 + z_tempyIntoNegCond1_G256_newbasis1);
    assign z6935_assgn6935 = dec_1_inp;
    assign z_x1_G256_newbasis1 = (t5 >> z2825_assgn2825);
    assign z_tempy2_G256_newbasis1 = z_y1_G256_newbasis1;
    assign z6941_assgn6941 = dec_1_inp;
    assign z_cond2_G256_newbasis1 = (z_x1_G256_newbasis1 & z2829_assgn2829);
    assign z_negCond2_G256_newbasis1 = !z_cond2_G256_newbasis1;
    assign z6947_assgn6947 = dec_3_inp;
    assign z_yxorb2_G256_newbasis1 = (z_y1_G256_newbasis1 ^ z2833_assgn2833);
    assign z_ny2_G256_newbasis1 = (z_cond2_G256_newbasis1 * z_yxorb2_G256_newbasis1);
    assign z_tempyIntoNegCond2_G256_newbasis1 = (z_tempy2_G256_newbasis1 * z_negCond2_G256_newbasis1);
    assign z_y2_G256_newbasis1 = (z_ny2_G256_newbasis1 + z_tempyIntoNegCond2_G256_newbasis1);
    assign z6957_assgn6957 = dec_1_inp;
    assign z_x2_G256_newbasis1 = (z_x1_G256_newbasis1 >> z2841_assgn2841);
    assign z_tempy3_G256_newbasis1 = z_y2_G256_newbasis1;
    assign z6963_assgn6963 = dec_1_inp;
    assign z_cond3_G256_newbasis1 = (z_x2_G256_newbasis1 & z2845_assgn2845);
    assign z_negCond3_G256_newbasis1 = !z_cond3_G256_newbasis1;
    assign z6969_assgn6969 = z3_assgn3;
    assign z_yxorb3_G256_newbasis1 = (z_y2_G256_newbasis1 ^ z2849_assgn2849);
    assign z_ny3_G256_newbasis1 = (z_cond3_G256_newbasis1 * z_yxorb3_G256_newbasis1);
    assign z_tempyIntoNegCond3_G256_newbasis1 = (z_tempy3_G256_newbasis1 * z_negCond3_G256_newbasis1);
    assign z_y3_G256_newbasis1 = (z_ny3_G256_newbasis1 + z_tempyIntoNegCond3_G256_newbasis1);
    assign z6979_assgn6979 = dec_1_inp;
    assign z_x3_G256_newbasis1 = (z_x2_G256_newbasis1 >> z2857_assgn2857);
    assign z_tempy4_G256_newbasis1 = z_y3_G256_newbasis1;
    assign z6985_assgn6985 = dec_1_inp;
    assign z_cond4_G256_newbasis1 = (z_x3_G256_newbasis1 & z2861_assgn2861);
    assign z_negCond4_G256_newbasis1 = !z_cond4_G256_newbasis1;
    assign z_yxorb4_G256_newbasis1 = (z_y3_G256_newbasis1 ^ dec_220_inp);
    assign z_ny4_G256_newbasis1 = (z_cond4_G256_newbasis1 * z_yxorb4_G256_newbasis1);
    assign z_tempyIntoNegCond4_G256_newbasis1 = (z_tempy4_G256_newbasis1 * z_negCond4_G256_newbasis1);
    assign z_y4_G256_newbasis1 = (z_ny4_G256_newbasis1 + z_tempyIntoNegCond4_G256_newbasis1);
    assign z6999_assgn6999 = dec_1_inp;
    assign z_x4_G256_newbasis1 = (z_x3_G256_newbasis1 >> z2873_assgn2873);
    assign z_tempy5_G256_newbasis1 = z_y4_G256_newbasis1;
    assign z7005_assgn7005 = dec_1_inp;
    assign z_cond5_G256_newbasis1 = (z_x4_G256_newbasis1 & z2877_assgn2877);
    assign z_negCond5_G256_newbasis1 = !z_cond5_G256_newbasis1;
    assign z_yxorb5_G256_newbasis1 = (z_y4_G256_newbasis1 ^ dec_11_inp);
    assign z_ny5_G256_newbasis1 = (z_cond5_G256_newbasis1 * z_yxorb5_G256_newbasis1);
    assign z_tempyIntoNegCond5_G256_newbasis1 = (z_tempy5_G256_newbasis1 * z_negCond5_G256_newbasis1);
    assign z_y5_G256_newbasis1 = (z_ny5_G256_newbasis1 + z_tempyIntoNegCond5_G256_newbasis1);
    assign z7019_assgn7019 = dec_1_inp;
    assign z_x5_G256_newbasis1 = (z_x4_G256_newbasis1 >> z2889_assgn2889);
    assign z_tempy6_G256_newbasis1 = z_y5_G256_newbasis1;
    assign z7025_assgn7025 = dec_1_inp;
    assign z_cond6_G256_newbasis1 = (z_x5_G256_newbasis1 & z2893_assgn2893);
    assign z_negCond6_G256_newbasis1 = !z_cond6_G256_newbasis1;
    assign z_yxorb6_G256_newbasis1 = (z_y5_G256_newbasis1 ^ dec_158_inp);
    assign z_ny6_G256_newbasis1 = (z_cond6_G256_newbasis1 * z_yxorb6_G256_newbasis1);
    assign z_tempyIntoNegCond6_G256_newbasis1 = (z_tempy6_G256_newbasis1 * z_negCond6_G256_newbasis1);
    assign z_y6_G256_newbasis1 = (z_ny6_G256_newbasis1 + z_tempyIntoNegCond6_G256_newbasis1);
    assign z7039_assgn7039 = dec_1_inp;
    assign z_x6_G256_newbasis1 = (z_x5_G256_newbasis1 >> z2905_assgn2905);
    assign z_tempy7_G256_newbasis1 = z_y6_G256_newbasis1;
    assign z7045_assgn7045 = dec_1_inp;
    assign z_cond7_G256_newbasis1 = (z_x6_G256_newbasis1 & z2909_assgn2909);
    assign z_negCond7_G256_newbasis1 = !z_cond7_G256_newbasis1;
    assign z_yxorb7_G256_newbasis1 = (z_y6_G256_newbasis1 ^ dec_45_inp);
    assign z_ny7_G256_newbasis1 = (z_cond7_G256_newbasis1 * z_yxorb7_G256_newbasis1);
    assign z_tempyIntoNegCond7_G256_newbasis1 = (z_tempy7_G256_newbasis1 * z_negCond7_G256_newbasis1);
    assign z_y7_G256_newbasis1 = (z_ny7_G256_newbasis1 + z_tempyIntoNegCond7_G256_newbasis1);
    assign z7059_assgn7059 = dec_1_inp;
    assign z_x7_G256_newbasis1 = (z_x6_G256_newbasis1 >> z2921_assgn2921);
    assign z_tempy8_G256_newbasis1 = z_y7_G256_newbasis1;
    assign z7065_assgn7065 = dec_1_inp;
    assign z_cond8_G256_newbasis1 = (z_x7_G256_newbasis1 & z2925_assgn2925);
    assign z_negCond8_G256_newbasis1 = !z_cond8_G256_newbasis1;
    assign z_yxorb8_G256_newbasis1 = (z_y7_G256_newbasis1 ^ dec_88_inp);
    assign z_ny8_G256_newbasis1 = (z_cond8_G256_newbasis1 * z_yxorb8_G256_newbasis1);
    assign z_tempyIntoNegCond8_G256_newbasis1 = (z_tempy8_G256_newbasis1 * z_negCond8_G256_newbasis1);
    assign z_y8_G256_newbasis1 = (z_ny8_G256_newbasis1 + z_tempyIntoNegCond8_G256_newbasis1);
    assign z7079_assgn7079 = dec_1_inp;
    assign z_x8_G256_newbasis1 = (z_x7_G256_newbasis1 >> z2937_assgn2937);
    assign t7 = z_y8_G256_newbasis1;

    always @(posedge clk) begin
        z2945_assgn29450 <= z2945_assgn2945;
        z2945_assgn29451 <= z2945_assgn29450;
        z2945_assgn29452 <= z2945_assgn29451;
        z2945_assgn29453 <= z2945_assgn29452;
        z2945_assgn29454 <= z2945_assgn29453;
        z2945_assgn29455 <= z2945_assgn29454;
        z2945_assgn29456 <= z2945_assgn29455;
        z2945_assgn29457 <= z2945_assgn29456;
        z2945_assgn29458 <= z2945_assgn29457;
        dec_99_inp <= z2945_assgn29458;
        z2947_assgn29470 <= z2947_assgn2947;
        z2947_assgn29471 <= z2947_assgn29470;
        z2947_assgn29472 <= z2947_assgn29471;
        z2947_assgn29473 <= z2947_assgn29472;
        z2947_assgn29474 <= z2947_assgn29473;
        z2947_assgn29475 <= z2947_assgn29474;
        z2947_assgn29476 <= z2947_assgn29475;
        z2947_assgn29477 <= z2947_assgn29476;
        z2947_assgn29478 <= z2947_assgn29477;
        dec_88_inp <= z2947_assgn29478;
        z2949_assgn29490 <= z2949_assgn2949;
        z2949_assgn29491 <= z2949_assgn29490;
        z2949_assgn29492 <= z2949_assgn29491;
        z2949_assgn29493 <= z2949_assgn29492;
        z2949_assgn29494 <= z2949_assgn29493;
        z2949_assgn29495 <= z2949_assgn29494;
        z2949_assgn29496 <= z2949_assgn29495;
        z2949_assgn29497 <= z2949_assgn29496;
        z2949_assgn29498 <= z2949_assgn29497;
        dec_45_inp <= z2949_assgn29498;
        z2951_assgn29510 <= z2951_assgn2951;
        z2951_assgn29511 <= z2951_assgn29510;
        z2951_assgn29512 <= z2951_assgn29511;
        z2951_assgn29513 <= z2951_assgn29512;
        z2951_assgn29514 <= z2951_assgn29513;
        z2951_assgn29515 <= z2951_assgn29514;
        z2951_assgn29516 <= z2951_assgn29515;
        z2951_assgn29517 <= z2951_assgn29516;
        z2951_assgn29518 <= z2951_assgn29517;
        dec_158_inp <= z2951_assgn29518;
        z2953_assgn29530 <= z2953_assgn2953;
        z2953_assgn29531 <= z2953_assgn29530;
        z2953_assgn29532 <= z2953_assgn29531;
        z2953_assgn29533 <= z2953_assgn29532;
        z2953_assgn29534 <= z2953_assgn29533;
        z2953_assgn29535 <= z2953_assgn29534;
        z2953_assgn29536 <= z2953_assgn29535;
        z2953_assgn29537 <= z2953_assgn29536;
        z2953_assgn29538 <= z2953_assgn29537;
        dec_11_inp <= z2953_assgn29538;
        z2955_assgn29550 <= z2955_assgn2955;
        z2955_assgn29551 <= z2955_assgn29550;
        z2955_assgn29552 <= z2955_assgn29551;
        z2955_assgn29553 <= z2955_assgn29552;
        z2955_assgn29554 <= z2955_assgn29553;
        z2955_assgn29555 <= z2955_assgn29554;
        z2955_assgn29556 <= z2955_assgn29555;
        z2955_assgn29557 <= z2955_assgn29556;
        z2955_assgn29558 <= z2955_assgn29557;
        dec_220_inp <= z2955_assgn29558;
        z2957_assgn29570 <= z2957_assgn2957;
        z2957_assgn29571 <= z2957_assgn29570;
        z2957_assgn29572 <= z2957_assgn29571;
        z2957_assgn29573 <= z2957_assgn29572;
        z2957_assgn29574 <= z2957_assgn29573;
        z2957_assgn29575 <= z2957_assgn29574;
        z2957_assgn29576 <= z2957_assgn29575;
        z2957_assgn29577 <= z2957_assgn29576;
        z2957_assgn29578 <= z2957_assgn29577;
        dec_36_inp <= z2957_assgn29578;
        z1_assgn1 <= dec_16_inp;
        z3_assgn3 <= dec_4_inp;
        z2975_assgn29750 <= z2975_assgn2975;
        z2975_assgn29751 <= z2975_assgn29750;
        dec_240_inp <= z2975_assgn29751;
        z5_assgn5 <= r0_inp;
        z7_assgn7 <= r1_inp;
        z9_assgn9 <= r2_inp;
        z11_assgn11 <= r3_inp;
        z13_assgn13 <= r4_inp;
        z15_assgn15 <= r5_inp;
        z17_assgn17 <= r6_inp;
        z19_assgn19 <= r7_inp;
        z21_assgn21 <= r8_inp;
        z3037_assgn30370 <= z3037_assgn3037;
        z3037_assgn30371 <= z3037_assgn30370;
        z3037_assgn30372 <= z3037_assgn30371;
        z3037_assgn30373 <= z3037_assgn30372;
        r9_inp <= z3037_assgn30373;
        z3039_assgn30390 <= z3039_assgn3039;
        z3039_assgn30391 <= z3039_assgn30390;
        z3039_assgn30392 <= z3039_assgn30391;
        z3039_assgn30393 <= z3039_assgn30392;
        r10_inp <= z3039_assgn30393;
        z3041_assgn30410 <= z3041_assgn3041;
        z3041_assgn30411 <= z3041_assgn30410;
        z3041_assgn30412 <= z3041_assgn30411;
        z3041_assgn30413 <= z3041_assgn30412;
        r11_inp <= z3041_assgn30413;
        z3043_assgn30430 <= z3043_assgn3043;
        z3043_assgn30431 <= z3043_assgn30430;
        z3043_assgn30432 <= z3043_assgn30431;
        z3043_assgn30433 <= z3043_assgn30432;
        z3043_assgn30434 <= z3043_assgn30433;
        r12_inp <= z3043_assgn30434;
        z3045_assgn30450 <= z3045_assgn3045;
        z3045_assgn30451 <= z3045_assgn30450;
        z3045_assgn30452 <= z3045_assgn30451;
        z3045_assgn30453 <= z3045_assgn30452;
        z3045_assgn30454 <= z3045_assgn30453;
        r13_inp <= z3045_assgn30454;
        z3047_assgn30470 <= z3047_assgn3047;
        z3047_assgn30471 <= z3047_assgn30470;
        z3047_assgn30472 <= z3047_assgn30471;
        z3047_assgn30473 <= z3047_assgn30472;
        z3047_assgn30474 <= z3047_assgn30473;
        r14_inp <= z3047_assgn30474;
        z3049_assgn30490 <= z3049_assgn3049;
        z3049_assgn30491 <= z3049_assgn30490;
        z3049_assgn30492 <= z3049_assgn30491;
        z3049_assgn30493 <= z3049_assgn30492;
        z3049_assgn30494 <= z3049_assgn30493;
        r15_inp <= z3049_assgn30494;
        z3051_assgn30510 <= z3051_assgn3051;
        z3051_assgn30511 <= z3051_assgn30510;
        z3051_assgn30512 <= z3051_assgn30511;
        z3051_assgn30513 <= z3051_assgn30512;
        z3051_assgn30514 <= z3051_assgn30513;
        r16_inp <= z3051_assgn30514;
        z3053_assgn30530 <= z3053_assgn3053;
        z3053_assgn30531 <= z3053_assgn30530;
        z3053_assgn30532 <= z3053_assgn30531;
        z3053_assgn30533 <= z3053_assgn30532;
        z3053_assgn30534 <= z3053_assgn30533;
        r17_inp <= z3053_assgn30534;
        z3055_assgn30550 <= z3055_assgn3055;
        z3055_assgn30551 <= z3055_assgn30550;
        z3055_assgn30552 <= z3055_assgn30551;
        z3055_assgn30553 <= z3055_assgn30552;
        z3055_assgn30554 <= z3055_assgn30553;
        z3055_assgn30555 <= z3055_assgn30554;
        r18_inp <= z3055_assgn30555;
        z3057_assgn30570 <= z3057_assgn3057;
        z3057_assgn30571 <= z3057_assgn30570;
        z3057_assgn30572 <= z3057_assgn30571;
        z3057_assgn30573 <= z3057_assgn30572;
        z3057_assgn30574 <= z3057_assgn30573;
        z3057_assgn30575 <= z3057_assgn30574;
        r19_inp <= z3057_assgn30575;
        z3059_assgn30590 <= z3059_assgn3059;
        z3059_assgn30591 <= z3059_assgn30590;
        z3059_assgn30592 <= z3059_assgn30591;
        z3059_assgn30593 <= z3059_assgn30592;
        z3059_assgn30594 <= z3059_assgn30593;
        z3059_assgn30595 <= z3059_assgn30594;
        r20_inp <= z3059_assgn30595;
        z3061_assgn30610 <= z3061_assgn3061;
        z3061_assgn30611 <= z3061_assgn30610;
        z3061_assgn30612 <= z3061_assgn30611;
        z3061_assgn30613 <= z3061_assgn30612;
        z3061_assgn30614 <= z3061_assgn30613;
        z3061_assgn30615 <= z3061_assgn30614;
        r21_inp <= z3061_assgn30615;
        z3063_assgn30630 <= z3063_assgn3063;
        z3063_assgn30631 <= z3063_assgn30630;
        z3063_assgn30632 <= z3063_assgn30631;
        z3063_assgn30633 <= z3063_assgn30632;
        z3063_assgn30634 <= z3063_assgn30633;
        z3063_assgn30635 <= z3063_assgn30634;
        r22_inp <= z3063_assgn30635;
        z3065_assgn30650 <= z3065_assgn3065;
        z3065_assgn30651 <= z3065_assgn30650;
        z3065_assgn30652 <= z3065_assgn30651;
        z3065_assgn30653 <= z3065_assgn30652;
        z3065_assgn30654 <= z3065_assgn30653;
        z3065_assgn30655 <= z3065_assgn30654;
        r23_inp <= z3065_assgn30655;
        z3067_assgn30670 <= z3067_assgn3067;
        z3067_assgn30671 <= z3067_assgn30670;
        z3067_assgn30672 <= z3067_assgn30671;
        z3067_assgn30673 <= z3067_assgn30672;
        z3067_assgn30674 <= z3067_assgn30673;
        z3067_assgn30675 <= z3067_assgn30674;
        r24_inp <= z3067_assgn30675;
        z3069_assgn30690 <= z3069_assgn3069;
        z3069_assgn30691 <= z3069_assgn30690;
        z3069_assgn30692 <= z3069_assgn30691;
        z3069_assgn30693 <= z3069_assgn30692;
        z3069_assgn30694 <= z3069_assgn30693;
        z3069_assgn30695 <= z3069_assgn30694;
        r25_inp <= z3069_assgn30695;
        z3071_assgn30710 <= z3071_assgn3071;
        z3071_assgn30711 <= z3071_assgn30710;
        z3071_assgn30712 <= z3071_assgn30711;
        z3071_assgn30713 <= z3071_assgn30712;
        z3071_assgn30714 <= z3071_assgn30713;
        z3071_assgn30715 <= z3071_assgn30714;
        r26_inp <= z3071_assgn30715;
        z3073_assgn30730 <= z3073_assgn3073;
        z3073_assgn30731 <= z3073_assgn30730;
        z3073_assgn30732 <= z3073_assgn30731;
        z3073_assgn30733 <= z3073_assgn30732;
        z3073_assgn30734 <= z3073_assgn30733;
        z3073_assgn30735 <= z3073_assgn30734;
        r27_inp <= z3073_assgn30735;
        z3075_assgn30750 <= z3075_assgn3075;
        z3075_assgn30751 <= z3075_assgn30750;
        z3075_assgn30752 <= z3075_assgn30751;
        z3075_assgn30753 <= z3075_assgn30752;
        z3075_assgn30754 <= z3075_assgn30753;
        z3075_assgn30755 <= z3075_assgn30754;
        r28_inp <= z3075_assgn30755;
        z3077_assgn30770 <= z3077_assgn3077;
        z3077_assgn30771 <= z3077_assgn30770;
        z3077_assgn30772 <= z3077_assgn30771;
        z3077_assgn30773 <= z3077_assgn30772;
        z3077_assgn30774 <= z3077_assgn30773;
        z3077_assgn30775 <= z3077_assgn30774;
        r29_inp <= z3077_assgn30775;
        z3079_assgn30790 <= z3079_assgn3079;
        z3079_assgn30791 <= z3079_assgn30790;
        z3079_assgn30792 <= z3079_assgn30791;
        z3079_assgn30793 <= z3079_assgn30792;
        z3079_assgn30794 <= z3079_assgn30793;
        z3079_assgn30795 <= z3079_assgn30794;
        r30_inp <= z3079_assgn30795;
        z3081_assgn30810 <= z3081_assgn3081;
        z3081_assgn30811 <= z3081_assgn30810;
        z3081_assgn30812 <= z3081_assgn30811;
        z3081_assgn30813 <= z3081_assgn30812;
        z3081_assgn30814 <= z3081_assgn30813;
        z3081_assgn30815 <= z3081_assgn30814;
        r31_inp <= z3081_assgn30815;
        z3083_assgn30830 <= z3083_assgn3083;
        z3083_assgn30831 <= z3083_assgn30830;
        z3083_assgn30832 <= z3083_assgn30831;
        z3083_assgn30833 <= z3083_assgn30832;
        z3083_assgn30834 <= z3083_assgn30833;
        z3083_assgn30835 <= z3083_assgn30834;
        r32_inp <= z3083_assgn30835;
        z3085_assgn30850 <= z3085_assgn3085;
        z3085_assgn30851 <= z3085_assgn30850;
        z3085_assgn30852 <= z3085_assgn30851;
        z3085_assgn30853 <= z3085_assgn30852;
        z3085_assgn30854 <= z3085_assgn30853;
        z3085_assgn30855 <= z3085_assgn30854;
        r33_inp <= z3085_assgn30855;
        z3087_assgn30870 <= z3087_assgn3087;
        z3087_assgn30871 <= z3087_assgn30870;
        z3087_assgn30872 <= z3087_assgn30871;
        z3087_assgn30873 <= z3087_assgn30872;
        z3087_assgn30874 <= z3087_assgn30873;
        z3087_assgn30875 <= z3087_assgn30874;
        r34_inp <= z3087_assgn30875;
        z3089_assgn30890 <= z3089_assgn3089;
        z3089_assgn30891 <= z3089_assgn30890;
        z3089_assgn30892 <= z3089_assgn30891;
        z3089_assgn30893 <= z3089_assgn30892;
        z3089_assgn30894 <= z3089_assgn30893;
        z3089_assgn30895 <= z3089_assgn30894;
        r35_inp <= z3089_assgn30895;
        z3219_assgn32190 <= z3219_assgn3219;
        z3219_assgn32191 <= z3219_assgn32190;
        z3219_assgn32192 <= z3219_assgn32191;
        z3219_assgn32193 <= z3219_assgn32192;
        z3219_assgn32194 <= z3219_assgn32193;
        z3219_assgn32195 <= z3219_assgn32194;
        z3219_assgn32196 <= z3219_assgn32195;
        z3219_assgn32197 <= z3219_assgn32196;
        z3219_assgn32198 <= z3219_assgn32197;
        z297_assgn297 <= z3219_assgn32198;
        z3221_assgn32210 <= z3221_assgn3221;
        z3221_assgn32211 <= z3221_assgn32210;
        z3221_assgn32212 <= z3221_assgn32211;
        z3221_assgn32213 <= z3221_assgn32212;
        z3221_assgn32214 <= z3221_assgn32213;
        z3221_assgn32215 <= z3221_assgn32214;
        z3221_assgn32216 <= z3221_assgn32215;
        z3221_assgn32217 <= z3221_assgn32216;
        z3221_assgn32218 <= z3221_assgn32217;
        z298_assgn298 <= z3221_assgn32218;
        z3355_assgn33550 <= z3355_assgn3355;
        z3355_assgn33551 <= z3355_assgn33550;
        z3355_assgn33552 <= z3355_assgn33551;
        z3355_assgn33553 <= z3355_assgn33552;
        z3355_assgn33554 <= z3355_assgn33553;
        z3355_assgn33555 <= z3355_assgn33554;
        z3355_assgn33556 <= z3355_assgn33555;
        z3355_assgn33557 <= z3355_assgn33556;
        z3355_assgn33558 <= z3355_assgn33557;
        z429_assgn429 <= z3355_assgn33558;
        z3357_assgn33570 <= z3357_assgn3357;
        z3357_assgn33571 <= z3357_assgn33570;
        z3357_assgn33572 <= z3357_assgn33571;
        z3357_assgn33573 <= z3357_assgn33572;
        z3357_assgn33574 <= z3357_assgn33573;
        z3357_assgn33575 <= z3357_assgn33574;
        z3357_assgn33576 <= z3357_assgn33575;
        z3357_assgn33577 <= z3357_assgn33576;
        z3357_assgn33578 <= z3357_assgn33577;
        z430_assgn430 <= z3357_assgn33578;
        z3363_assgn33630 <= z3363_assgn3363;
        z3363_assgn33631 <= z3363_assgn33630;
        z434_assgn434 <= z3363_assgn33631;
        z3367_assgn33670 <= z3367_assgn3367;
        z3367_assgn33671 <= z3367_assgn33670;
        z436_assgn436 <= z3367_assgn33671;
        z3371_assgn33710 <= z3371_assgn3371;
        z437_assgn437 <= z3371_assgn33710;
        z3375_assgn33750 <= z3375_assgn3375;
        z439_assgn439 <= z3375_assgn33750;
        z3383_assgn33830 <= z3383_assgn3383;
        z3383_assgn33831 <= z3383_assgn33830;
        z3383_assgn33832 <= z3383_assgn33831;
        z445_assgn445 <= z3383_assgn33832;
        a0_G256_inv0_reg <= a0_G256_inv0;
        z3387_assgn33870 <= z3387_assgn3387;
        z3387_assgn33871 <= z3387_assgn33870;
        z3387_assgn33872 <= z3387_assgn33871;
        z447_assgn447 <= z3387_assgn33872;
        a1_G256_inv0_reg <= a1_G256_inv0;
        z3391_assgn33910 <= z3391_assgn3391;
        z3391_assgn33911 <= z3391_assgn33910;
        z3391_assgn33912 <= z3391_assgn33911;
        z449_assgn449 <= z3391_assgn33912;
        z3395_assgn33950 <= z3395_assgn3395;
        z3395_assgn33951 <= z3395_assgn33950;
        z3395_assgn33952 <= z3395_assgn33951;
        z451_assgn451 <= z3395_assgn33952;
        z3399_assgn33990 <= z3399_assgn3399;
        z3399_assgn33991 <= z3399_assgn33990;
        z3399_assgn33992 <= z3399_assgn33991;
        z453_assgn453 <= z3399_assgn33992;
        z3403_assgn34030 <= z3403_assgn3403;
        z3403_assgn34031 <= z3403_assgn34030;
        z3403_assgn34032 <= z3403_assgn34031;
        z455_assgn455 <= z3403_assgn34032;
        z3407_assgn34070 <= z3407_assgn3407;
        z3407_assgn34071 <= z3407_assgn34070;
        z3407_assgn34072 <= z3407_assgn34071;
        z457_assgn457 <= z3407_assgn34072;
        z3411_assgn34110 <= z3411_assgn3411;
        z3411_assgn34111 <= z3411_assgn34110;
        z3411_assgn34112 <= z3411_assgn34111;
        z459_assgn459 <= z3411_assgn34112;
        z3419_assgn34190 <= z3419_assgn3419;
        z3419_assgn34191 <= z3419_assgn34190;
        z3419_assgn34192 <= z3419_assgn34191;
        z465_assgn465 <= z3419_assgn34192;
        z3423_assgn34230 <= z3423_assgn3423;
        z3423_assgn34231 <= z3423_assgn34230;
        z3423_assgn34232 <= z3423_assgn34231;
        z467_assgn467 <= z3423_assgn34232;
        z3427_assgn34270 <= z3427_assgn3427;
        z3427_assgn34271 <= z3427_assgn34270;
        z3427_assgn34272 <= z3427_assgn34271;
        z469_assgn469 <= z3427_assgn34272;
        z3431_assgn34310 <= z3431_assgn3431;
        z3431_assgn34311 <= z3431_assgn34310;
        z3431_assgn34312 <= z3431_assgn34311;
        z471_assgn471 <= z3431_assgn34312;
        z3435_assgn34350 <= z3435_assgn3435;
        z3435_assgn34351 <= z3435_assgn34350;
        z3435_assgn34352 <= z3435_assgn34351;
        z473_assgn473 <= z3435_assgn34352;
        z3439_assgn34390 <= z3439_assgn3439;
        z3439_assgn34391 <= z3439_assgn34390;
        z3439_assgn34392 <= z3439_assgn34391;
        z475_assgn475 <= z3439_assgn34392;
        z3443_assgn34430 <= z3443_assgn3443;
        z3443_assgn34431 <= z3443_assgn34430;
        z3443_assgn34432 <= z3443_assgn34431;
        z477_assgn477 <= z3443_assgn34432;
        z3447_assgn34470 <= z3447_assgn3447;
        z3447_assgn34471 <= z3447_assgn34470;
        z3447_assgn34472 <= z3447_assgn34471;
        z479_assgn479 <= z3447_assgn34472;
        z3455_assgn34550 <= z3455_assgn3455;
        z3455_assgn34551 <= z3455_assgn34550;
        z3455_assgn34552 <= z3455_assgn34551;
        z485_assgn485 <= z3455_assgn34552;
        z3459_assgn34590 <= z3459_assgn3459;
        z3459_assgn34591 <= z3459_assgn34590;
        z3459_assgn34592 <= z3459_assgn34591;
        z487_assgn487 <= z3459_assgn34592;
        z3463_assgn34630 <= z3463_assgn3463;
        z3463_assgn34631 <= z3463_assgn34630;
        z3463_assgn34632 <= z3463_assgn34631;
        z489_assgn489 <= z3463_assgn34632;
        z3467_assgn34670 <= z3467_assgn3467;
        z3467_assgn34671 <= z3467_assgn34670;
        z3467_assgn34672 <= z3467_assgn34671;
        z491_assgn491 <= z3467_assgn34672;
        z3471_assgn34710 <= z3471_assgn3471;
        z3471_assgn34711 <= z3471_assgn34710;
        z3471_assgn34712 <= z3471_assgn34711;
        z493_assgn493 <= z3471_assgn34712;
        z3475_assgn34750 <= z3475_assgn3475;
        z3475_assgn34751 <= z3475_assgn34750;
        z3475_assgn34752 <= z3475_assgn34751;
        z495_assgn495 <= z3475_assgn34752;
        z3479_assgn34790 <= z3479_assgn3479;
        z3479_assgn34791 <= z3479_assgn34790;
        z3479_assgn34792 <= z3479_assgn34791;
        z497_assgn497 <= z3479_assgn34792;
        z3483_assgn34830 <= z3483_assgn3483;
        z3483_assgn34831 <= z3483_assgn34830;
        z3483_assgn34832 <= z3483_assgn34831;
        z499_assgn499 <= z3483_assgn34832;
        z3491_assgn34910 <= z3491_assgn3491;
        z3491_assgn34911 <= z3491_assgn34910;
        z3491_assgn34912 <= z3491_assgn34911;
        z505_assgn505 <= z3491_assgn34912;
        z3495_assgn34950 <= z3495_assgn3495;
        z3495_assgn34951 <= z3495_assgn34950;
        z3495_assgn34952 <= z3495_assgn34951;
        z507_assgn507 <= z3495_assgn34952;
        z3499_assgn34990 <= z3499_assgn3499;
        z3499_assgn34991 <= z3499_assgn34990;
        z3499_assgn34992 <= z3499_assgn34991;
        z509_assgn509 <= z3499_assgn34992;
        z3503_assgn35030 <= z3503_assgn3503;
        z3503_assgn35031 <= z3503_assgn35030;
        z3503_assgn35032 <= z3503_assgn35031;
        z511_assgn511 <= z3503_assgn35032;
        z3507_assgn35070 <= z3507_assgn3507;
        z3507_assgn35071 <= z3507_assgn35070;
        z3507_assgn35072 <= z3507_assgn35071;
        z513_assgn513 <= z3507_assgn35072;
        z3511_assgn35110 <= z3511_assgn3511;
        z3511_assgn35111 <= z3511_assgn35110;
        z3511_assgn35112 <= z3511_assgn35111;
        z515_assgn515 <= z3511_assgn35112;
        z3523_assgn35230 <= z3523_assgn3523;
        z3523_assgn35231 <= z3523_assgn35230;
        z3523_assgn35232 <= z3523_assgn35231;
        z525_assgn525 <= z3523_assgn35232;
        z3527_assgn35270 <= z3527_assgn3527;
        z3527_assgn35271 <= z3527_assgn35270;
        z3527_assgn35272 <= z3527_assgn35271;
        z527_assgn527 <= z3527_assgn35272;
        z3535_assgn35350 <= z3535_assgn3535;
        z3535_assgn35351 <= z3535_assgn35350;
        z3535_assgn35352 <= z3535_assgn35351;
        z533_assgn533 <= z3535_assgn35352;
        z3539_assgn35390 <= z3539_assgn3539;
        z3539_assgn35391 <= z3539_assgn35390;
        z3539_assgn35392 <= z3539_assgn35391;
        z535_assgn535 <= z3539_assgn35392;
        z3565_assgn35650 <= z3565_assgn3565;
        z3565_assgn35651 <= z3565_assgn35650;
        z559_assgn559 <= z3565_assgn35651;
        z3569_assgn35690 <= z3569_assgn3569;
        z3569_assgn35691 <= z3569_assgn35690;
        z561_assgn561 <= z3569_assgn35691;
        z3573_assgn35730 <= z3573_assgn3573;
        z3573_assgn35731 <= z3573_assgn35730;
        z563_assgn563 <= z3573_assgn35731;
        z3577_assgn35770 <= z3577_assgn3577;
        z3577_assgn35771 <= z3577_assgn35770;
        z565_assgn565 <= z3577_assgn35771;
        z3581_assgn35810 <= z3581_assgn3581;
        z3581_assgn35811 <= z3581_assgn35810;
        z567_assgn567 <= z3581_assgn35811;
        z3585_assgn35850 <= z3585_assgn3585;
        z3585_assgn35851 <= z3585_assgn35850;
        z569_assgn569 <= z3585_assgn35851;
        z3615_assgn36150 <= z3615_assgn3615;
        z3615_assgn36151 <= z3615_assgn36150;
        z597_assgn597 <= z3615_assgn36151;
        z3619_assgn36190 <= z3619_assgn3619;
        z3619_assgn36191 <= z3619_assgn36190;
        z599_assgn599 <= z3619_assgn36191;
        z3623_assgn36230 <= z3623_assgn3623;
        z3623_assgn36231 <= z3623_assgn36230;
        z601_assgn601 <= z3623_assgn36231;
        z3627_assgn36270 <= z3627_assgn3627;
        z3627_assgn36271 <= z3627_assgn36270;
        z603_assgn603 <= z3627_assgn36271;
        z3631_assgn36310 <= z3631_assgn3631;
        z3631_assgn36311 <= z3631_assgn36310;
        z605_assgn605 <= z3631_assgn36311;
        z3635_assgn36350 <= z3635_assgn3635;
        z3635_assgn36351 <= z3635_assgn36350;
        z607_assgn607 <= z3635_assgn36351;
        c0_G4_mul0_G16_mul0_G256_inv0_reg <= c0_G4_mul0_G16_mul0_G256_inv0;
        d0_G4_mul0_G16_mul0_G256_inv0_reg <= d0_G4_mul0_G16_mul0_G256_inv0;
        c1_G4_mul0_G16_mul0_G256_inv0_reg <= c1_G4_mul0_G16_mul0_G256_inv0;
        d1_G4_mul0_G16_mul0_G256_inv0_reg <= d1_G4_mul0_G16_mul0_G256_inv0;
        dec_2_inp_reg <= dec_2_inp;
        z3665_assgn36650 <= z3665_assgn3665;
        z635_assgn635 <= z3665_assgn36650;
        z3669_assgn36690 <= z3669_assgn3669;
        z637_assgn637 <= z3669_assgn36690;
        cxord_0_G4_mul0_G16_mul0_G256_inv0_reg <= cxord_0_G4_mul0_G16_mul0_G256_inv0;
        r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= r0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        cxord_1_G4_mul0_G16_mul0_G256_inv0_reg <= cxord_1_G4_mul0_G16_mul0_G256_inv0;
        z3677_assgn36770 <= z3677_assgn3677;
        z643_assgn643 <= z3677_assgn36770;
        v1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= v1_hpc20_G4_mul0_G16_mul0_G256_inv0;
        u0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= u0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        z3687_assgn36870 <= z3687_assgn3687;
        z651_assgn651 <= z3687_assgn36870;
        v0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= v0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        u1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= u1_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p3_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p3_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p2_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p2_hpc20_G4_mul0_G16_mul0_G256_inv0;
        z3703_assgn37030 <= z3703_assgn3703;
        z665_assgn665 <= z3703_assgn37030;
        z3707_assgn37070 <= z3707_assgn3707;
        z667_assgn667 <= z3707_assgn37070;
        z3711_assgn37110 <= z3711_assgn3711;
        z670_assgn670 <= z3711_assgn37110;
        r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= r0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        z3715_assgn37150 <= z3715_assgn3715;
        z672_assgn672 <= z3715_assgn37150;
        z3719_assgn37190 <= z3719_assgn3719;
        z3719_assgn37191 <= z3719_assgn37190;
        z673_assgn673 <= z3719_assgn37191;
        v1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= v1_hpc21_G4_mul0_G16_mul0_G256_inv0;
        u0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= u0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        z3729_assgn37290 <= z3729_assgn3729;
        z3729_assgn37291 <= z3729_assgn37290;
        z681_assgn681 <= z3729_assgn37291;
        v0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= v0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        u1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= u1_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p3_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p3_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p2_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p2_hpc21_G4_mul0_G16_mul0_G256_inv0;
        z3749_assgn37490 <= z3749_assgn3749;
        z699_assgn699 <= z3749_assgn37490;
        z3753_assgn37530 <= z3753_assgn3753;
        z701_assgn701 <= z3753_assgn37530;
        z3757_assgn37570 <= z3757_assgn3757;
        z704_assgn704 <= z3757_assgn37570;
        r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= r0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        z3761_assgn37610 <= z3761_assgn3761;
        z706_assgn706 <= z3761_assgn37610;
        z3765_assgn37650 <= z3765_assgn3765;
        z3765_assgn37651 <= z3765_assgn37650;
        z707_assgn707 <= z3765_assgn37651;
        v1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= v1_hpc22_G4_mul0_G16_mul0_G256_inv0;
        u0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= u0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        z3775_assgn37750 <= z3775_assgn3775;
        z3775_assgn37751 <= z3775_assgn37750;
        z715_assgn715 <= z3775_assgn37751;
        v0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= v0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        u1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= u1_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p3_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p3_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p2_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p2_hpc22_G4_mul0_G16_mul0_G256_inv0;
        z3789_assgn37890 <= z3789_assgn3789;
        z3789_assgn37891 <= z3789_assgn37890;
        z3789_assgn37892 <= z3789_assgn37891;
        z727_assgn727 <= z3789_assgn37892;
        z3793_assgn37930 <= z3793_assgn3793;
        z3793_assgn37931 <= z3793_assgn37930;
        z3793_assgn37932 <= z3793_assgn37931;
        z729_assgn729 <= z3793_assgn37932;
        z3801_assgn38010 <= z3801_assgn3801;
        z3801_assgn38011 <= z3801_assgn38010;
        z3801_assgn38012 <= z3801_assgn38011;
        z735_assgn735 <= z3801_assgn38012;
        z3805_assgn38050 <= z3805_assgn3805;
        z3805_assgn38051 <= z3805_assgn38050;
        z3805_assgn38052 <= z3805_assgn38051;
        z737_assgn737 <= z3805_assgn38052;
        z3809_assgn38090 <= z3809_assgn3809;
        z3809_assgn38091 <= z3809_assgn38090;
        z3809_assgn38092 <= z3809_assgn38091;
        z739_assgn739 <= z3809_assgn38092;
        z3813_assgn38130 <= z3813_assgn3813;
        z3813_assgn38131 <= z3813_assgn38130;
        z3813_assgn38132 <= z3813_assgn38131;
        z741_assgn741 <= z3813_assgn38132;
        z3817_assgn38170 <= z3817_assgn3817;
        z3817_assgn38171 <= z3817_assgn38170;
        z3817_assgn38172 <= z3817_assgn38171;
        z743_assgn743 <= z3817_assgn38172;
        z3821_assgn38210 <= z3821_assgn3821;
        z3821_assgn38211 <= z3821_assgn38210;
        z3821_assgn38212 <= z3821_assgn38211;
        z745_assgn745 <= z3821_assgn38212;
        z3833_assgn38330 <= z3833_assgn3833;
        z3833_assgn38331 <= z3833_assgn38330;
        z3833_assgn38332 <= z3833_assgn38331;
        z755_assgn755 <= z3833_assgn38332;
        z3837_assgn38370 <= z3837_assgn3837;
        z3837_assgn38371 <= z3837_assgn38370;
        z3837_assgn38372 <= z3837_assgn38371;
        z757_assgn757 <= z3837_assgn38372;
        z3851_assgn38510 <= z3851_assgn3851;
        z3851_assgn38511 <= z3851_assgn38510;
        z769_assgn769 <= z3851_assgn38511;
        z3855_assgn38550 <= z3855_assgn3855;
        z3855_assgn38551 <= z3855_assgn38550;
        z771_assgn771 <= z3855_assgn38551;
        z3859_assgn38590 <= z3859_assgn3859;
        z3859_assgn38591 <= z3859_assgn38590;
        z773_assgn773 <= z3859_assgn38591;
        z3863_assgn38630 <= z3863_assgn3863;
        z3863_assgn38631 <= z3863_assgn38630;
        z775_assgn775 <= z3863_assgn38631;
        z3867_assgn38670 <= z3867_assgn3867;
        z3867_assgn38671 <= z3867_assgn38670;
        z777_assgn777 <= z3867_assgn38671;
        z3871_assgn38710 <= z3871_assgn3871;
        z3871_assgn38711 <= z3871_assgn38710;
        z779_assgn779 <= z3871_assgn38711;
        c0_G4_mul1_G16_mul0_G256_inv0_reg <= c0_G4_mul1_G16_mul0_G256_inv0;
        d0_G4_mul1_G16_mul0_G256_inv0_reg <= d0_G4_mul1_G16_mul0_G256_inv0;
        c1_G4_mul1_G16_mul0_G256_inv0_reg <= c1_G4_mul1_G16_mul0_G256_inv0;
        d1_G4_mul1_G16_mul0_G256_inv0_reg <= d1_G4_mul1_G16_mul0_G256_inv0;
        z3901_assgn39010 <= z3901_assgn3901;
        z807_assgn807 <= z3901_assgn39010;
        z3905_assgn39050 <= z3905_assgn3905;
        z809_assgn809 <= z3905_assgn39050;
        cxord_0_G4_mul1_G16_mul0_G256_inv0_reg <= cxord_0_G4_mul1_G16_mul0_G256_inv0;
        r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= r0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        cxord_1_G4_mul1_G16_mul0_G256_inv0_reg <= cxord_1_G4_mul1_G16_mul0_G256_inv0;
        z3913_assgn39130 <= z3913_assgn3913;
        z815_assgn815 <= z3913_assgn39130;
        v1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= v1_hpc20_G4_mul1_G16_mul0_G256_inv0;
        u0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= u0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        z3923_assgn39230 <= z3923_assgn3923;
        z823_assgn823 <= z3923_assgn39230;
        v0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= v0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        u1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= u1_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p3_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p3_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p2_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p2_hpc20_G4_mul1_G16_mul0_G256_inv0;
        z3939_assgn39390 <= z3939_assgn3939;
        z837_assgn837 <= z3939_assgn39390;
        z3943_assgn39430 <= z3943_assgn3943;
        z839_assgn839 <= z3943_assgn39430;
        z3947_assgn39470 <= z3947_assgn3947;
        z842_assgn842 <= z3947_assgn39470;
        r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= r0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        z3951_assgn39510 <= z3951_assgn3951;
        z844_assgn844 <= z3951_assgn39510;
        z3955_assgn39550 <= z3955_assgn3955;
        z3955_assgn39551 <= z3955_assgn39550;
        z845_assgn845 <= z3955_assgn39551;
        v1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= v1_hpc21_G4_mul1_G16_mul0_G256_inv0;
        u0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= u0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        z3965_assgn39650 <= z3965_assgn3965;
        z3965_assgn39651 <= z3965_assgn39650;
        z853_assgn853 <= z3965_assgn39651;
        v0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= v0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        u1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= u1_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p3_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p3_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p2_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p2_hpc21_G4_mul1_G16_mul0_G256_inv0;
        z3985_assgn39850 <= z3985_assgn3985;
        z871_assgn871 <= z3985_assgn39850;
        z3989_assgn39890 <= z3989_assgn3989;
        z873_assgn873 <= z3989_assgn39890;
        z3993_assgn39930 <= z3993_assgn3993;
        z876_assgn876 <= z3993_assgn39930;
        r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= r0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        z3997_assgn39970 <= z3997_assgn3997;
        z878_assgn878 <= z3997_assgn39970;
        z4001_assgn40010 <= z4001_assgn4001;
        z4001_assgn40011 <= z4001_assgn40010;
        z879_assgn879 <= z4001_assgn40011;
        v1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= v1_hpc22_G4_mul1_G16_mul0_G256_inv0;
        u0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= u0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        z4011_assgn40110 <= z4011_assgn4011;
        z4011_assgn40111 <= z4011_assgn40110;
        z887_assgn887 <= z4011_assgn40111;
        v0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= v0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        u1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= u1_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p3_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p3_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p2_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p2_hpc22_G4_mul1_G16_mul0_G256_inv0;
        z4025_assgn40250 <= z4025_assgn4025;
        z4025_assgn40251 <= z4025_assgn40250;
        z4025_assgn40252 <= z4025_assgn40251;
        z899_assgn899 <= z4025_assgn40252;
        z4029_assgn40290 <= z4029_assgn4029;
        z4029_assgn40291 <= z4029_assgn40290;
        z4029_assgn40292 <= z4029_assgn40291;
        z901_assgn901 <= z4029_assgn40292;
        z4047_assgn40470 <= z4047_assgn4047;
        z4047_assgn40471 <= z4047_assgn40470;
        z917_assgn917 <= z4047_assgn40471;
        z4051_assgn40510 <= z4051_assgn4051;
        z4051_assgn40511 <= z4051_assgn40510;
        z919_assgn919 <= z4051_assgn40511;
        z4055_assgn40550 <= z4055_assgn4055;
        z4055_assgn40551 <= z4055_assgn40550;
        z921_assgn921 <= z4055_assgn40551;
        z4059_assgn40590 <= z4059_assgn4059;
        z4059_assgn40591 <= z4059_assgn40590;
        z923_assgn923 <= z4059_assgn40591;
        z4063_assgn40630 <= z4063_assgn4063;
        z4063_assgn40631 <= z4063_assgn40630;
        z925_assgn925 <= z4063_assgn40631;
        z4067_assgn40670 <= z4067_assgn4067;
        z4067_assgn40671 <= z4067_assgn40670;
        z927_assgn927 <= z4067_assgn40671;
        c0_G4_mul2_G16_mul0_G256_inv0_reg <= c0_G4_mul2_G16_mul0_G256_inv0;
        d0_G4_mul2_G16_mul0_G256_inv0_reg <= d0_G4_mul2_G16_mul0_G256_inv0;
        c1_G4_mul2_G16_mul0_G256_inv0_reg <= c1_G4_mul2_G16_mul0_G256_inv0;
        d1_G4_mul2_G16_mul0_G256_inv0_reg <= d1_G4_mul2_G16_mul0_G256_inv0;
        z4097_assgn40970 <= z4097_assgn4097;
        z955_assgn955 <= z4097_assgn40970;
        z4101_assgn41010 <= z4101_assgn4101;
        z957_assgn957 <= z4101_assgn41010;
        cxord_0_G4_mul2_G16_mul0_G256_inv0_reg <= cxord_0_G4_mul2_G16_mul0_G256_inv0;
        r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= r0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        cxord_1_G4_mul2_G16_mul0_G256_inv0_reg <= cxord_1_G4_mul2_G16_mul0_G256_inv0;
        z4109_assgn41090 <= z4109_assgn4109;
        z963_assgn963 <= z4109_assgn41090;
        v1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= v1_hpc20_G4_mul2_G16_mul0_G256_inv0;
        u0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= u0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        z4119_assgn41190 <= z4119_assgn4119;
        z971_assgn971 <= z4119_assgn41190;
        v0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= v0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        u1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= u1_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p3_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p3_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p2_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p2_hpc20_G4_mul2_G16_mul0_G256_inv0;
        z4135_assgn41350 <= z4135_assgn4135;
        z985_assgn985 <= z4135_assgn41350;
        z4139_assgn41390 <= z4139_assgn4139;
        z987_assgn987 <= z4139_assgn41390;
        z4143_assgn41430 <= z4143_assgn4143;
        z990_assgn990 <= z4143_assgn41430;
        r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= r0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        z4147_assgn41470 <= z4147_assgn4147;
        z992_assgn992 <= z4147_assgn41470;
        z4151_assgn41510 <= z4151_assgn4151;
        z4151_assgn41511 <= z4151_assgn41510;
        z993_assgn993 <= z4151_assgn41511;
        v1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= v1_hpc21_G4_mul2_G16_mul0_G256_inv0;
        u0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= u0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        z4161_assgn41610 <= z4161_assgn4161;
        z4161_assgn41611 <= z4161_assgn41610;
        z1001_assgn1001 <= z4161_assgn41611;
        v0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= v0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        u1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= u1_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p3_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p3_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p2_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p2_hpc21_G4_mul2_G16_mul0_G256_inv0;
        z4181_assgn41810 <= z4181_assgn4181;
        z1019_assgn1019 <= z4181_assgn41810;
        z4185_assgn41850 <= z4185_assgn4185;
        z1021_assgn1021 <= z4185_assgn41850;
        z4189_assgn41890 <= z4189_assgn4189;
        z1024_assgn1024 <= z4189_assgn41890;
        r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= r0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        z4193_assgn41930 <= z4193_assgn4193;
        z1026_assgn1026 <= z4193_assgn41930;
        z4197_assgn41970 <= z4197_assgn4197;
        z4197_assgn41971 <= z4197_assgn41970;
        z1027_assgn1027 <= z4197_assgn41971;
        v1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= v1_hpc22_G4_mul2_G16_mul0_G256_inv0;
        u0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= u0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        z4207_assgn42070 <= z4207_assgn4207;
        z4207_assgn42071 <= z4207_assgn42070;
        z1035_assgn1035 <= z4207_assgn42071;
        v0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= v0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        u1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= u1_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p3_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p3_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p2_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p2_hpc22_G4_mul2_G16_mul0_G256_inv0;
        z4221_assgn42210 <= z4221_assgn4221;
        z4221_assgn42211 <= z4221_assgn42210;
        z4221_assgn42212 <= z4221_assgn42211;
        z1047_assgn1047 <= z4221_assgn42212;
        z4225_assgn42250 <= z4225_assgn4225;
        z4225_assgn42251 <= z4225_assgn42250;
        z4225_assgn42252 <= z4225_assgn42251;
        z1049_assgn1049 <= z4225_assgn42252;
        z4237_assgn42370 <= z4237_assgn4237;
        z4237_assgn42371 <= z4237_assgn42370;
        z4237_assgn42372 <= z4237_assgn42371;
        z1059_assgn1059 <= z4237_assgn42372;
        z4241_assgn42410 <= z4241_assgn4241;
        z4241_assgn42411 <= z4241_assgn42410;
        z4241_assgn42412 <= z4241_assgn42411;
        z1061_assgn1061 <= z4241_assgn42412;
        z4253_assgn42530 <= z4253_assgn4253;
        z4253_assgn42531 <= z4253_assgn42530;
        z4253_assgn42532 <= z4253_assgn42531;
        z1071_assgn1071 <= z4253_assgn42532;
        z4257_assgn42570 <= z4257_assgn4257;
        z4257_assgn42571 <= z4257_assgn42570;
        z4257_assgn42572 <= z4257_assgn42571;
        z1073_assgn1073 <= z4257_assgn42572;
        z4261_assgn42610 <= z4261_assgn4261;
        z4261_assgn42611 <= z4261_assgn42610;
        z4261_assgn42612 <= z4261_assgn42611;
        z1075_assgn1075 <= z4261_assgn42612;
        z4265_assgn42650 <= z4265_assgn4265;
        z4265_assgn42651 <= z4265_assgn42650;
        z4265_assgn42652 <= z4265_assgn42651;
        z4265_assgn42653 <= z4265_assgn42652;
        z1077_assgn1077 <= z4265_assgn42653;
        z4269_assgn42690 <= z4269_assgn4269;
        z4269_assgn42691 <= z4269_assgn42690;
        z4269_assgn42692 <= z4269_assgn42691;
        z4269_assgn42693 <= z4269_assgn42692;
        z1079_assgn1079 <= z4269_assgn42693;
        z4273_assgn42730 <= z4273_assgn4273;
        z4273_assgn42731 <= z4273_assgn42730;
        z4273_assgn42732 <= z4273_assgn42731;
        z4273_assgn42733 <= z4273_assgn42732;
        z1081_assgn1081 <= z4273_assgn42733;
        z4277_assgn42770 <= z4277_assgn4277;
        z4277_assgn42771 <= z4277_assgn42770;
        z4277_assgn42772 <= z4277_assgn42771;
        z4277_assgn42773 <= z4277_assgn42772;
        z1083_assgn1083 <= z4277_assgn42773;
        z4281_assgn42810 <= z4281_assgn4281;
        z4281_assgn42811 <= z4281_assgn42810;
        z4281_assgn42812 <= z4281_assgn42811;
        z4281_assgn42813 <= z4281_assgn42812;
        z1085_assgn1085 <= z4281_assgn42813;
        z4285_assgn42850 <= z4285_assgn4285;
        z4285_assgn42851 <= z4285_assgn42850;
        z4285_assgn42852 <= z4285_assgn42851;
        z4285_assgn42853 <= z4285_assgn42852;
        z1087_assgn1087 <= z4285_assgn42853;
        z4289_assgn42890 <= z4289_assgn4289;
        z4289_assgn42891 <= z4289_assgn42890;
        z4289_assgn42892 <= z4289_assgn42891;
        z4289_assgn42893 <= z4289_assgn42892;
        z1089_assgn1089 <= z4289_assgn42893;
        c0xord0_G256_inv0_reg <= c0xord0_G256_inv0;
        z4293_assgn42930 <= z4293_assgn4293;
        z4293_assgn42931 <= z4293_assgn42930;
        z4293_assgn42932 <= z4293_assgn42931;
        z4293_assgn42933 <= z4293_assgn42932;
        z1091_assgn1091 <= z4293_assgn42933;
        c1xord1_G256_inv0_reg <= c1xord1_G256_inv0;
        z4297_assgn42970 <= z4297_assgn4297;
        z4297_assgn42971 <= z4297_assgn42970;
        z4297_assgn42972 <= z4297_assgn42971;
        z4297_assgn42973 <= z4297_assgn42972;
        z1093_assgn1093 <= z4297_assgn42973;
        z4301_assgn43010 <= z4301_assgn4301;
        z4301_assgn43011 <= z4301_assgn43010;
        z4301_assgn43012 <= z4301_assgn43011;
        z4301_assgn43013 <= z4301_assgn43012;
        z1095_assgn1095 <= z4301_assgn43013;
        z4305_assgn43050 <= z4305_assgn4305;
        z4305_assgn43051 <= z4305_assgn43050;
        z4305_assgn43052 <= z4305_assgn43051;
        z1097_assgn1097 <= z4305_assgn43052;
        z4309_assgn43090 <= z4309_assgn4309;
        z4309_assgn43091 <= z4309_assgn43090;
        z4309_assgn43092 <= z4309_assgn43091;
        z1099_assgn1099 <= z4309_assgn43092;
        z4313_assgn43130 <= z4313_assgn4313;
        z4313_assgn43131 <= z4313_assgn43130;
        z4313_assgn43132 <= z4313_assgn43131;
        z1101_assgn1101 <= z4313_assgn43132;
        z4315_assgn43150 <= z4315_assgn4315;
        z4315_assgn43151 <= z4315_assgn43150;
        z1102_assgn1102 <= z4315_assgn43151;
        z4319_assgn43190 <= z4319_assgn4319;
        z4319_assgn43191 <= z4319_assgn43190;
        z4319_assgn43192 <= z4319_assgn43191;
        z1103_assgn1103 <= z4319_assgn43192;
        z4321_assgn43210 <= z4321_assgn4321;
        z4321_assgn43211 <= z4321_assgn43210;
        z1104_assgn1104 <= z4321_assgn43211;
        z4325_assgn43250 <= z4325_assgn4325;
        z4325_assgn43251 <= z4325_assgn43250;
        z4325_assgn43252 <= z4325_assgn43251;
        z4325_assgn43253 <= z4325_assgn43252;
        z4325_assgn43254 <= z4325_assgn43253;
        z4325_assgn43255 <= z4325_assgn43254;
        z4325_assgn43256 <= z4325_assgn43255;
        z1105_assgn1105 <= z4325_assgn43256;
        z4329_assgn43290 <= z4329_assgn4329;
        z4329_assgn43291 <= z4329_assgn43290;
        z4329_assgn43292 <= z4329_assgn43291;
        z4329_assgn43293 <= z4329_assgn43292;
        z4329_assgn43294 <= z4329_assgn43293;
        z4329_assgn43295 <= z4329_assgn43294;
        z4329_assgn43296 <= z4329_assgn43295;
        z1107_assgn1107 <= z4329_assgn43296;
        z4333_assgn43330 <= z4333_assgn4333;
        z4333_assgn43331 <= z4333_assgn43330;
        z4333_assgn43332 <= z4333_assgn43331;
        z4333_assgn43333 <= z4333_assgn43332;
        z4333_assgn43334 <= z4333_assgn43333;
        z4333_assgn43335 <= z4333_assgn43334;
        z4333_assgn43336 <= z4333_assgn43335;
        z1109_assgn1109 <= z4333_assgn43336;
        z4337_assgn43370 <= z4337_assgn4337;
        z4337_assgn43371 <= z4337_assgn43370;
        z4337_assgn43372 <= z4337_assgn43371;
        z4337_assgn43373 <= z4337_assgn43372;
        z4337_assgn43374 <= z4337_assgn43373;
        z4337_assgn43375 <= z4337_assgn43374;
        z4337_assgn43376 <= z4337_assgn43375;
        z1111_assgn1111 <= z4337_assgn43376;
        z4341_assgn43410 <= z4341_assgn4341;
        z4341_assgn43411 <= z4341_assgn43410;
        z4341_assgn43412 <= z4341_assgn43411;
        z4341_assgn43413 <= z4341_assgn43412;
        z4341_assgn43414 <= z4341_assgn43413;
        z4341_assgn43415 <= z4341_assgn43414;
        z4341_assgn43416 <= z4341_assgn43415;
        z1113_assgn1113 <= z4341_assgn43416;
        z4345_assgn43450 <= z4345_assgn4345;
        z4345_assgn43451 <= z4345_assgn43450;
        z4345_assgn43452 <= z4345_assgn43451;
        z4345_assgn43453 <= z4345_assgn43452;
        z4345_assgn43454 <= z4345_assgn43453;
        z4345_assgn43455 <= z4345_assgn43454;
        z4345_assgn43456 <= z4345_assgn43455;
        z1115_assgn1115 <= z4345_assgn43456;
        z4349_assgn43490 <= z4349_assgn4349;
        z4349_assgn43491 <= z4349_assgn43490;
        z4349_assgn43492 <= z4349_assgn43491;
        z4349_assgn43493 <= z4349_assgn43492;
        z4349_assgn43494 <= z4349_assgn43493;
        z4349_assgn43495 <= z4349_assgn43494;
        z4349_assgn43496 <= z4349_assgn43495;
        z1117_assgn1117 <= z4349_assgn43496;
        z4353_assgn43530 <= z4353_assgn4353;
        z4353_assgn43531 <= z4353_assgn43530;
        z4353_assgn43532 <= z4353_assgn43531;
        z4353_assgn43533 <= z4353_assgn43532;
        z4353_assgn43534 <= z4353_assgn43533;
        z4353_assgn43535 <= z4353_assgn43534;
        z4353_assgn43536 <= z4353_assgn43535;
        z1119_assgn1119 <= z4353_assgn43536;
        z4361_assgn43610 <= z4361_assgn4361;
        z4361_assgn43611 <= z4361_assgn43610;
        z4361_assgn43612 <= z4361_assgn43611;
        z4361_assgn43613 <= z4361_assgn43612;
        z4361_assgn43614 <= z4361_assgn43613;
        z4361_assgn43615 <= z4361_assgn43614;
        z4361_assgn43616 <= z4361_assgn43615;
        z1125_assgn1125 <= z4361_assgn43616;
        z4365_assgn43650 <= z4365_assgn4365;
        z4365_assgn43651 <= z4365_assgn43650;
        z4365_assgn43652 <= z4365_assgn43651;
        z4365_assgn43653 <= z4365_assgn43652;
        z4365_assgn43654 <= z4365_assgn43653;
        z4365_assgn43655 <= z4365_assgn43654;
        z4365_assgn43656 <= z4365_assgn43655;
        z1127_assgn1127 <= z4365_assgn43656;
        z4369_assgn43690 <= z4369_assgn4369;
        z4369_assgn43691 <= z4369_assgn43690;
        z4369_assgn43692 <= z4369_assgn43691;
        z4369_assgn43693 <= z4369_assgn43692;
        z4369_assgn43694 <= z4369_assgn43693;
        z4369_assgn43695 <= z4369_assgn43694;
        z4369_assgn43696 <= z4369_assgn43695;
        z1129_assgn1129 <= z4369_assgn43696;
        z4373_assgn43730 <= z4373_assgn4373;
        z4373_assgn43731 <= z4373_assgn43730;
        z4373_assgn43732 <= z4373_assgn43731;
        z4373_assgn43733 <= z4373_assgn43732;
        z4373_assgn43734 <= z4373_assgn43733;
        z4373_assgn43735 <= z4373_assgn43734;
        z4373_assgn43736 <= z4373_assgn43735;
        z1131_assgn1131 <= z4373_assgn43736;
        z4377_assgn43770 <= z4377_assgn4377;
        z4377_assgn43771 <= z4377_assgn43770;
        z4377_assgn43772 <= z4377_assgn43771;
        z4377_assgn43773 <= z4377_assgn43772;
        z4377_assgn43774 <= z4377_assgn43773;
        z4377_assgn43775 <= z4377_assgn43774;
        z4377_assgn43776 <= z4377_assgn43775;
        z1133_assgn1133 <= z4377_assgn43776;
        z4381_assgn43810 <= z4381_assgn4381;
        z4381_assgn43811 <= z4381_assgn43810;
        z4381_assgn43812 <= z4381_assgn43811;
        z4381_assgn43813 <= z4381_assgn43812;
        z4381_assgn43814 <= z4381_assgn43813;
        z4381_assgn43815 <= z4381_assgn43814;
        z4381_assgn43816 <= z4381_assgn43815;
        z1135_assgn1135 <= z4381_assgn43816;
        z4393_assgn43930 <= z4393_assgn4393;
        z4393_assgn43931 <= z4393_assgn43930;
        z4393_assgn43932 <= z4393_assgn43931;
        z4393_assgn43933 <= z4393_assgn43932;
        z4393_assgn43934 <= z4393_assgn43933;
        z4393_assgn43935 <= z4393_assgn43934;
        z4393_assgn43936 <= z4393_assgn43935;
        z1145_assgn1145 <= z4393_assgn43936;
        z4397_assgn43970 <= z4397_assgn4397;
        z4397_assgn43971 <= z4397_assgn43970;
        z4397_assgn43972 <= z4397_assgn43971;
        z4397_assgn43973 <= z4397_assgn43972;
        z4397_assgn43974 <= z4397_assgn43973;
        z4397_assgn43975 <= z4397_assgn43974;
        z4397_assgn43976 <= z4397_assgn43975;
        z1147_assgn1147 <= z4397_assgn43976;
        z4405_assgn44050 <= z4405_assgn4405;
        z4405_assgn44051 <= z4405_assgn44050;
        z4405_assgn44052 <= z4405_assgn44051;
        z1153_assgn1153 <= z4405_assgn44052;
        z4409_assgn44090 <= z4409_assgn4409;
        z4409_assgn44091 <= z4409_assgn44090;
        z4409_assgn44092 <= z4409_assgn44091;
        z1155_assgn1155 <= z4409_assgn44092;
        z4413_assgn44130 <= z4413_assgn4413;
        z4413_assgn44131 <= z4413_assgn44130;
        z4413_assgn44132 <= z4413_assgn44131;
        z1157_assgn1157 <= z4413_assgn44132;
        z4417_assgn44170 <= z4417_assgn4417;
        z4417_assgn44171 <= z4417_assgn44170;
        z4417_assgn44172 <= z4417_assgn44171;
        z4417_assgn44173 <= z4417_assgn44172;
        z4417_assgn44174 <= z4417_assgn44173;
        z4417_assgn44175 <= z4417_assgn44174;
        z1159_assgn1159 <= z4417_assgn44175;
        z4419_assgn44190 <= z4419_assgn4419;
        z1160_assgn1160 <= z4419_assgn44190;
        z4423_assgn44230 <= z4423_assgn4423;
        z4423_assgn44231 <= z4423_assgn44230;
        z4423_assgn44232 <= z4423_assgn44231;
        z4423_assgn44233 <= z4423_assgn44232;
        z4423_assgn44234 <= z4423_assgn44233;
        z4423_assgn44235 <= z4423_assgn44234;
        z1161_assgn1161 <= z4423_assgn44235;
        z4425_assgn44250 <= z4425_assgn4425;
        z1162_assgn1162 <= z4425_assgn44250;
        z4429_assgn44290 <= z4429_assgn4429;
        z4429_assgn44291 <= z4429_assgn44290;
        z4429_assgn44292 <= z4429_assgn44291;
        z4429_assgn44293 <= z4429_assgn44292;
        z4429_assgn44294 <= z4429_assgn44293;
        z4429_assgn44295 <= z4429_assgn44294;
        z1163_assgn1163 <= z4429_assgn44295;
        z4433_assgn44330 <= z4433_assgn4433;
        z4433_assgn44331 <= z4433_assgn44330;
        z4433_assgn44332 <= z4433_assgn44331;
        z4433_assgn44333 <= z4433_assgn44332;
        z4433_assgn44334 <= z4433_assgn44333;
        z4433_assgn44335 <= z4433_assgn44334;
        z1165_assgn1165 <= z4433_assgn44335;
        z4437_assgn44370 <= z4437_assgn4437;
        z4437_assgn44371 <= z4437_assgn44370;
        z4437_assgn44372 <= z4437_assgn44371;
        z4437_assgn44373 <= z4437_assgn44372;
        z4437_assgn44374 <= z4437_assgn44373;
        z4437_assgn44375 <= z4437_assgn44374;
        z1167_assgn1167 <= z4437_assgn44375;
        z4439_assgn44390 <= z4439_assgn4439;
        z1168_assgn1168 <= z4439_assgn44390;
        z4443_assgn44430 <= z4443_assgn4443;
        z4443_assgn44431 <= z4443_assgn44430;
        z4443_assgn44432 <= z4443_assgn44431;
        z4443_assgn44433 <= z4443_assgn44432;
        z4443_assgn44434 <= z4443_assgn44433;
        z4443_assgn44435 <= z4443_assgn44434;
        z1169_assgn1169 <= z4443_assgn44435;
        z4445_assgn44450 <= z4445_assgn4445;
        z1170_assgn1170 <= z4445_assgn44450;
        z4449_assgn44490 <= z4449_assgn4449;
        z4449_assgn44491 <= z4449_assgn44490;
        z4449_assgn44492 <= z4449_assgn44491;
        z1171_assgn1171 <= z4449_assgn44492;
        z4453_assgn44530 <= z4453_assgn4453;
        z4453_assgn44531 <= z4453_assgn44530;
        z4453_assgn44532 <= z4453_assgn44531;
        z1173_assgn1173 <= z4453_assgn44532;
        z4457_assgn44570 <= z4457_assgn4457;
        z4457_assgn44571 <= z4457_assgn44570;
        z4457_assgn44572 <= z4457_assgn44571;
        z1175_assgn1175 <= z4457_assgn44572;
        z4461_assgn44610 <= z4461_assgn4461;
        z4461_assgn44611 <= z4461_assgn44610;
        z4461_assgn44612 <= z4461_assgn44611;
        z1177_assgn1177 <= z4461_assgn44612;
        z4465_assgn44650 <= z4465_assgn4465;
        z4465_assgn44651 <= z4465_assgn44650;
        z4465_assgn44652 <= z4465_assgn44651;
        z1179_assgn1179 <= z4465_assgn44652;
        z4469_assgn44690 <= z4469_assgn4469;
        z4469_assgn44691 <= z4469_assgn44690;
        z4469_assgn44692 <= z4469_assgn44691;
        z1181_assgn1181 <= z4469_assgn44692;
        c0_G4_mul3_G16_inv0_G256_inv0_reg <= c0_G4_mul3_G16_inv0_G256_inv0;
        d0_G4_mul3_G16_inv0_G256_inv0_reg <= d0_G4_mul3_G16_inv0_G256_inv0;
        c1_G4_mul3_G16_inv0_G256_inv0_reg <= c1_G4_mul3_G16_inv0_G256_inv0;
        d1_G4_mul3_G16_inv0_G256_inv0_reg <= d1_G4_mul3_G16_inv0_G256_inv0;
        z4481_assgn44810 <= z4481_assgn4481;
        z4481_assgn44811 <= z4481_assgn44810;
        z4481_assgn44812 <= z4481_assgn44811;
        z4481_assgn44813 <= z4481_assgn44812;
        z1191_assgn1191 <= z4481_assgn44813;
        z4489_assgn44890 <= z4489_assgn4489;
        z1197_assgn1197 <= z4489_assgn44890;
        z4493_assgn44930 <= z4493_assgn4493;
        z1199_assgn1199 <= z4493_assgn44930;
        cxord_0_G4_mul3_G16_inv0_G256_inv0_reg <= cxord_0_G4_mul3_G16_inv0_G256_inv0;
        r0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
        cxord_1_G4_mul3_G16_inv0_G256_inv0_reg <= cxord_1_G4_mul3_G16_inv0_G256_inv0;
        z4501_assgn45010 <= z4501_assgn4501;
        z1205_assgn1205 <= z4501_assgn45010;
        v1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= v1_hpc20_G4_mul3_G16_inv0_G256_inv0;
        u0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= u0_hpc20_G4_mul3_G16_inv0_G256_inv0;
        p1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc20_G4_mul3_G16_inv0_G256_inv0;
        p0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p0_hpc20_G4_mul3_G16_inv0_G256_inv0;
        z4511_assgn45110 <= z4511_assgn4511;
        z1213_assgn1213 <= z4511_assgn45110;
        v0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= v0_hpc20_G4_mul3_G16_inv0_G256_inv0;
        u1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= u1_hpc20_G4_mul3_G16_inv0_G256_inv0;
        p3_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p3_hpc20_G4_mul3_G16_inv0_G256_inv0;
        p2_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p2_hpc20_G4_mul3_G16_inv0_G256_inv0;
        z4521_assgn45210 <= z4521_assgn4521;
        z4521_assgn45211 <= z4521_assgn45210;
        z4521_assgn45212 <= z4521_assgn45211;
        z4521_assgn45213 <= z4521_assgn45212;
        z1221_assgn1221 <= z4521_assgn45213;
        z4529_assgn45290 <= z4529_assgn4529;
        z1227_assgn1227 <= z4529_assgn45290;
        z4533_assgn45330 <= z4533_assgn4533;
        z1229_assgn1229 <= z4533_assgn45330;
        z4537_assgn45370 <= z4537_assgn4537;
        z1232_assgn1232 <= z4537_assgn45370;
        r0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
        z4541_assgn45410 <= z4541_assgn4541;
        z1234_assgn1234 <= z4541_assgn45410;
        z4545_assgn45450 <= z4545_assgn4545;
        z4545_assgn45451 <= z4545_assgn45450;
        z1235_assgn1235 <= z4545_assgn45451;
        v1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= v1_hpc21_G4_mul3_G16_inv0_G256_inv0;
        u0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= u0_hpc21_G4_mul3_G16_inv0_G256_inv0;
        p1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc21_G4_mul3_G16_inv0_G256_inv0;
        p0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p0_hpc21_G4_mul3_G16_inv0_G256_inv0;
        z4555_assgn45550 <= z4555_assgn4555;
        z4555_assgn45551 <= z4555_assgn45550;
        z1243_assgn1243 <= z4555_assgn45551;
        v0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= v0_hpc21_G4_mul3_G16_inv0_G256_inv0;
        u1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= u1_hpc21_G4_mul3_G16_inv0_G256_inv0;
        p3_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p3_hpc21_G4_mul3_G16_inv0_G256_inv0;
        p2_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p2_hpc21_G4_mul3_G16_inv0_G256_inv0;
        z4569_assgn45690 <= z4569_assgn4569;
        z4569_assgn45691 <= z4569_assgn45690;
        z4569_assgn45692 <= z4569_assgn45691;
        z4569_assgn45693 <= z4569_assgn45692;
        z1255_assgn1255 <= z4569_assgn45693;
        z4577_assgn45770 <= z4577_assgn4577;
        z1261_assgn1261 <= z4577_assgn45770;
        z4581_assgn45810 <= z4581_assgn4581;
        z1263_assgn1263 <= z4581_assgn45810;
        z4585_assgn45850 <= z4585_assgn4585;
        z1266_assgn1266 <= z4585_assgn45850;
        r0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
        z4589_assgn45890 <= z4589_assgn4589;
        z1268_assgn1268 <= z4589_assgn45890;
        z4593_assgn45930 <= z4593_assgn4593;
        z4593_assgn45931 <= z4593_assgn45930;
        z1269_assgn1269 <= z4593_assgn45931;
        v1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= v1_hpc22_G4_mul3_G16_inv0_G256_inv0;
        u0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= u0_hpc22_G4_mul3_G16_inv0_G256_inv0;
        p1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc22_G4_mul3_G16_inv0_G256_inv0;
        p0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p0_hpc22_G4_mul3_G16_inv0_G256_inv0;
        z4603_assgn46030 <= z4603_assgn4603;
        z4603_assgn46031 <= z4603_assgn46030;
        z1277_assgn1277 <= z4603_assgn46031;
        v0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= v0_hpc22_G4_mul3_G16_inv0_G256_inv0;
        u1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= u1_hpc22_G4_mul3_G16_inv0_G256_inv0;
        p3_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p3_hpc22_G4_mul3_G16_inv0_G256_inv0;
        p2_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p2_hpc22_G4_mul3_G16_inv0_G256_inv0;
        z4617_assgn46170 <= z4617_assgn4617;
        z4617_assgn46171 <= z4617_assgn46170;
        z4617_assgn46172 <= z4617_assgn46171;
        z4617_assgn46173 <= z4617_assgn46172;
        z4617_assgn46174 <= z4617_assgn46173;
        z4617_assgn46175 <= z4617_assgn46174;
        z4617_assgn46176 <= z4617_assgn46175;
        z1289_assgn1289 <= z4617_assgn46176;
        z4621_assgn46210 <= z4621_assgn4621;
        z4621_assgn46211 <= z4621_assgn46210;
        z4621_assgn46212 <= z4621_assgn46211;
        z4621_assgn46213 <= z4621_assgn46212;
        z4621_assgn46214 <= z4621_assgn46213;
        z4621_assgn46215 <= z4621_assgn46214;
        z4621_assgn46216 <= z4621_assgn46215;
        z1291_assgn1291 <= z4621_assgn46216;
        z4633_assgn46330 <= z4633_assgn4633;
        z4633_assgn46331 <= z4633_assgn46330;
        z4633_assgn46332 <= z4633_assgn46331;
        z4633_assgn46333 <= z4633_assgn46332;
        z4633_assgn46334 <= z4633_assgn46333;
        z4633_assgn46335 <= z4633_assgn46334;
        z4633_assgn46336 <= z4633_assgn46335;
        z1301_assgn1301 <= z4633_assgn46336;
        z4637_assgn46370 <= z4637_assgn4637;
        z4637_assgn46371 <= z4637_assgn46370;
        z4637_assgn46372 <= z4637_assgn46371;
        z4637_assgn46373 <= z4637_assgn46372;
        z4637_assgn46374 <= z4637_assgn46373;
        z4637_assgn46375 <= z4637_assgn46374;
        z4637_assgn46376 <= z4637_assgn46375;
        z1303_assgn1303 <= z4637_assgn46376;
        z4641_assgn46410 <= z4641_assgn4641;
        z4641_assgn46411 <= z4641_assgn46410;
        z4641_assgn46412 <= z4641_assgn46411;
        z4641_assgn46413 <= z4641_assgn46412;
        z4641_assgn46414 <= z4641_assgn46413;
        z4641_assgn46415 <= z4641_assgn46414;
        z4641_assgn46416 <= z4641_assgn46415;
        z1305_assgn1305 <= z4641_assgn46416;
        z4645_assgn46450 <= z4645_assgn4645;
        z4645_assgn46451 <= z4645_assgn46450;
        z4645_assgn46452 <= z4645_assgn46451;
        z4645_assgn46453 <= z4645_assgn46452;
        z4645_assgn46454 <= z4645_assgn46453;
        z4645_assgn46455 <= z4645_assgn46454;
        z4645_assgn46456 <= z4645_assgn46455;
        z1307_assgn1307 <= z4645_assgn46456;
        z4649_assgn46490 <= z4649_assgn4649;
        z4649_assgn46491 <= z4649_assgn46490;
        z4649_assgn46492 <= z4649_assgn46491;
        z4649_assgn46493 <= z4649_assgn46492;
        z4649_assgn46494 <= z4649_assgn46493;
        z4649_assgn46495 <= z4649_assgn46494;
        z4649_assgn46496 <= z4649_assgn46495;
        z1309_assgn1309 <= z4649_assgn46496;
        z4653_assgn46530 <= z4653_assgn4653;
        z4653_assgn46531 <= z4653_assgn46530;
        z4653_assgn46532 <= z4653_assgn46531;
        z4653_assgn46533 <= z4653_assgn46532;
        z4653_assgn46534 <= z4653_assgn46533;
        z4653_assgn46535 <= z4653_assgn46534;
        z4653_assgn46536 <= z4653_assgn46535;
        z1311_assgn1311 <= z4653_assgn46536;
        z4657_assgn46570 <= z4657_assgn4657;
        z4657_assgn46571 <= z4657_assgn46570;
        z4657_assgn46572 <= z4657_assgn46571;
        z4657_assgn46573 <= z4657_assgn46572;
        z4657_assgn46574 <= z4657_assgn46573;
        z4657_assgn46575 <= z4657_assgn46574;
        z4657_assgn46576 <= z4657_assgn46575;
        z1313_assgn1313 <= z4657_assgn46576;
        z4661_assgn46610 <= z4661_assgn4661;
        z4661_assgn46611 <= z4661_assgn46610;
        z4661_assgn46612 <= z4661_assgn46611;
        z4661_assgn46613 <= z4661_assgn46612;
        z4661_assgn46614 <= z4661_assgn46613;
        z4661_assgn46615 <= z4661_assgn46614;
        z4661_assgn46616 <= z4661_assgn46615;
        z1315_assgn1315 <= z4661_assgn46616;
        z4669_assgn46690 <= z4669_assgn4669;
        z4669_assgn46691 <= z4669_assgn46690;
        z4669_assgn46692 <= z4669_assgn46691;
        z4669_assgn46693 <= z4669_assgn46692;
        z1321_assgn1321 <= z4669_assgn46693;
        z4673_assgn46730 <= z4673_assgn4673;
        z4673_assgn46731 <= z4673_assgn46730;
        z4673_assgn46732 <= z4673_assgn46731;
        z4673_assgn46733 <= z4673_assgn46732;
        z1323_assgn1323 <= z4673_assgn46733;
        z4677_assgn46770 <= z4677_assgn4677;
        z4677_assgn46771 <= z4677_assgn46770;
        z4677_assgn46772 <= z4677_assgn46771;
        z4677_assgn46773 <= z4677_assgn46772;
        z1325_assgn1325 <= z4677_assgn46773;
        z4681_assgn46810 <= z4681_assgn4681;
        z4681_assgn46811 <= z4681_assgn46810;
        z4681_assgn46812 <= z4681_assgn46811;
        z4681_assgn46813 <= z4681_assgn46812;
        z4681_assgn46814 <= z4681_assgn46813;
        z4681_assgn46815 <= z4681_assgn46814;
        z4681_assgn46816 <= z4681_assgn46815;
        z1327_assgn1327 <= z4681_assgn46816;
        z4685_assgn46850 <= z4685_assgn4685;
        z4685_assgn46851 <= z4685_assgn46850;
        z4685_assgn46852 <= z4685_assgn46851;
        z4685_assgn46853 <= z4685_assgn46852;
        z4685_assgn46854 <= z4685_assgn46853;
        z4685_assgn46855 <= z4685_assgn46854;
        z4685_assgn46856 <= z4685_assgn46855;
        z1329_assgn1329 <= z4685_assgn46856;
        z4689_assgn46890 <= z4689_assgn4689;
        z4689_assgn46891 <= z4689_assgn46890;
        z4689_assgn46892 <= z4689_assgn46891;
        z4689_assgn46893 <= z4689_assgn46892;
        z4689_assgn46894 <= z4689_assgn46893;
        z4689_assgn46895 <= z4689_assgn46894;
        z4689_assgn46896 <= z4689_assgn46895;
        z1331_assgn1331 <= z4689_assgn46896;
        z4693_assgn46930 <= z4693_assgn4693;
        z4693_assgn46931 <= z4693_assgn46930;
        z4693_assgn46932 <= z4693_assgn46931;
        z4693_assgn46933 <= z4693_assgn46932;
        z4693_assgn46934 <= z4693_assgn46933;
        z4693_assgn46935 <= z4693_assgn46934;
        z4693_assgn46936 <= z4693_assgn46935;
        z1333_assgn1333 <= z4693_assgn46936;
        z4697_assgn46970 <= z4697_assgn4697;
        z4697_assgn46971 <= z4697_assgn46970;
        z4697_assgn46972 <= z4697_assgn46971;
        z4697_assgn46973 <= z4697_assgn46972;
        z4697_assgn46974 <= z4697_assgn46973;
        z4697_assgn46975 <= z4697_assgn46974;
        z4697_assgn46976 <= z4697_assgn46975;
        z1335_assgn1335 <= z4697_assgn46976;
        z4701_assgn47010 <= z4701_assgn4701;
        z4701_assgn47011 <= z4701_assgn47010;
        z4701_assgn47012 <= z4701_assgn47011;
        z4701_assgn47013 <= z4701_assgn47012;
        z4701_assgn47014 <= z4701_assgn47013;
        z4701_assgn47015 <= z4701_assgn47014;
        z4701_assgn47016 <= z4701_assgn47015;
        z1337_assgn1337 <= z4701_assgn47016;
        z4705_assgn47050 <= z4705_assgn4705;
        z4705_assgn47051 <= z4705_assgn47050;
        z4705_assgn47052 <= z4705_assgn47051;
        z4705_assgn47053 <= z4705_assgn47052;
        z1339_assgn1339 <= z4705_assgn47053;
        b0_G16_inv0_G256_inv0_reg <= b0_G16_inv0_G256_inv0;
        z4709_assgn47090 <= z4709_assgn4709;
        z4709_assgn47091 <= z4709_assgn47090;
        z4709_assgn47092 <= z4709_assgn47091;
        z4709_assgn47093 <= z4709_assgn47092;
        z1341_assgn1341 <= z4709_assgn47093;
        b1_G16_inv0_G256_inv0_reg <= b1_G16_inv0_G256_inv0;
        z4713_assgn47130 <= z4713_assgn4713;
        z4713_assgn47131 <= z4713_assgn47130;
        z4713_assgn47132 <= z4713_assgn47131;
        z4713_assgn47133 <= z4713_assgn47132;
        z1343_assgn1343 <= z4713_assgn47133;
        z4717_assgn47170 <= z4717_assgn4717;
        z4717_assgn47171 <= z4717_assgn47170;
        z4717_assgn47172 <= z4717_assgn47171;
        z4717_assgn47173 <= z4717_assgn47172;
        z1345_assgn1345 <= z4717_assgn47173;
        z4721_assgn47210 <= z4721_assgn4721;
        z4721_assgn47211 <= z4721_assgn47210;
        z4721_assgn47212 <= z4721_assgn47211;
        z4721_assgn47213 <= z4721_assgn47212;
        z1347_assgn1347 <= z4721_assgn47213;
        z4725_assgn47250 <= z4725_assgn4725;
        z4725_assgn47251 <= z4725_assgn47250;
        z4725_assgn47252 <= z4725_assgn47251;
        z4725_assgn47253 <= z4725_assgn47252;
        z1349_assgn1349 <= z4725_assgn47253;
        c0_G4_mul4_G16_inv0_G256_inv0_reg <= c0_G4_mul4_G16_inv0_G256_inv0;
        d0_G4_mul4_G16_inv0_G256_inv0_reg <= d0_G4_mul4_G16_inv0_G256_inv0;
        c1_G4_mul4_G16_inv0_G256_inv0_reg <= c1_G4_mul4_G16_inv0_G256_inv0;
        d1_G4_mul4_G16_inv0_G256_inv0_reg <= d1_G4_mul4_G16_inv0_G256_inv0;
        z4737_assgn47370 <= z4737_assgn4737;
        z4737_assgn47371 <= z4737_assgn47370;
        z4737_assgn47372 <= z4737_assgn47371;
        z4737_assgn47373 <= z4737_assgn47372;
        z4737_assgn47374 <= z4737_assgn47373;
        z1359_assgn1359 <= z4737_assgn47374;
        z4745_assgn47450 <= z4745_assgn4745;
        z1365_assgn1365 <= z4745_assgn47450;
        z4749_assgn47490 <= z4749_assgn4749;
        z1367_assgn1367 <= z4749_assgn47490;
        cxord_0_G4_mul4_G16_inv0_G256_inv0_reg <= cxord_0_G4_mul4_G16_inv0_G256_inv0;
        r0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
        cxord_1_G4_mul4_G16_inv0_G256_inv0_reg <= cxord_1_G4_mul4_G16_inv0_G256_inv0;
        z4757_assgn47570 <= z4757_assgn4757;
        z1373_assgn1373 <= z4757_assgn47570;
        v1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= v1_hpc20_G4_mul4_G16_inv0_G256_inv0;
        u0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= u0_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p0_hpc20_G4_mul4_G16_inv0_G256_inv0;
        z4767_assgn47670 <= z4767_assgn4767;
        z1381_assgn1381 <= z4767_assgn47670;
        v0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= v0_hpc20_G4_mul4_G16_inv0_G256_inv0;
        u1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= u1_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p3_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p3_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p2_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p2_hpc20_G4_mul4_G16_inv0_G256_inv0;
        z4777_assgn47770 <= z4777_assgn4777;
        z4777_assgn47771 <= z4777_assgn47770;
        z4777_assgn47772 <= z4777_assgn47771;
        z4777_assgn47773 <= z4777_assgn47772;
        z4777_assgn47774 <= z4777_assgn47773;
        z1389_assgn1389 <= z4777_assgn47774;
        z4785_assgn47850 <= z4785_assgn4785;
        z1395_assgn1395 <= z4785_assgn47850;
        z4789_assgn47890 <= z4789_assgn4789;
        z1397_assgn1397 <= z4789_assgn47890;
        z4793_assgn47930 <= z4793_assgn4793;
        z1400_assgn1400 <= z4793_assgn47930;
        r0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
        z4797_assgn47970 <= z4797_assgn4797;
        z1402_assgn1402 <= z4797_assgn47970;
        z4801_assgn48010 <= z4801_assgn4801;
        z4801_assgn48011 <= z4801_assgn48010;
        z1403_assgn1403 <= z4801_assgn48011;
        v1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= v1_hpc21_G4_mul4_G16_inv0_G256_inv0;
        u0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= u0_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p0_hpc21_G4_mul4_G16_inv0_G256_inv0;
        z4811_assgn48110 <= z4811_assgn4811;
        z4811_assgn48111 <= z4811_assgn48110;
        z1411_assgn1411 <= z4811_assgn48111;
        v0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= v0_hpc21_G4_mul4_G16_inv0_G256_inv0;
        u1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= u1_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p3_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p3_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p2_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p2_hpc21_G4_mul4_G16_inv0_G256_inv0;
        z4825_assgn48250 <= z4825_assgn4825;
        z4825_assgn48251 <= z4825_assgn48250;
        z4825_assgn48252 <= z4825_assgn48251;
        z4825_assgn48253 <= z4825_assgn48252;
        z4825_assgn48254 <= z4825_assgn48253;
        z1423_assgn1423 <= z4825_assgn48254;
        z4833_assgn48330 <= z4833_assgn4833;
        z1429_assgn1429 <= z4833_assgn48330;
        z4837_assgn48370 <= z4837_assgn4837;
        z1431_assgn1431 <= z4837_assgn48370;
        z4841_assgn48410 <= z4841_assgn4841;
        z1434_assgn1434 <= z4841_assgn48410;
        r0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
        z4845_assgn48450 <= z4845_assgn4845;
        z1436_assgn1436 <= z4845_assgn48450;
        z4849_assgn48490 <= z4849_assgn4849;
        z4849_assgn48491 <= z4849_assgn48490;
        z1437_assgn1437 <= z4849_assgn48491;
        v1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= v1_hpc22_G4_mul4_G16_inv0_G256_inv0;
        u0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= u0_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p0_hpc22_G4_mul4_G16_inv0_G256_inv0;
        z4859_assgn48590 <= z4859_assgn4859;
        z4859_assgn48591 <= z4859_assgn48590;
        z1445_assgn1445 <= z4859_assgn48591;
        v0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= v0_hpc22_G4_mul4_G16_inv0_G256_inv0;
        u1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= u1_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p3_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p3_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p2_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p2_hpc22_G4_mul4_G16_inv0_G256_inv0;
        z4873_assgn48730 <= z4873_assgn4873;
        z4873_assgn48731 <= z4873_assgn48730;
        z4873_assgn48732 <= z4873_assgn48731;
        z4873_assgn48733 <= z4873_assgn48732;
        z4873_assgn48734 <= z4873_assgn48733;
        z4873_assgn48735 <= z4873_assgn48734;
        z4873_assgn48736 <= z4873_assgn48735;
        z4873_assgn48737 <= z4873_assgn48736;
        z1457_assgn1457 <= z4873_assgn48737;
        z4877_assgn48770 <= z4877_assgn4877;
        z4877_assgn48771 <= z4877_assgn48770;
        z4877_assgn48772 <= z4877_assgn48771;
        z4877_assgn48773 <= z4877_assgn48772;
        z4877_assgn48774 <= z4877_assgn48773;
        z4877_assgn48775 <= z4877_assgn48774;
        z4877_assgn48776 <= z4877_assgn48775;
        z4877_assgn48777 <= z4877_assgn48776;
        z1459_assgn1459 <= z4877_assgn48777;
        z4885_assgn48850 <= z4885_assgn4885;
        z4885_assgn48851 <= z4885_assgn48850;
        z4885_assgn48852 <= z4885_assgn48851;
        z4885_assgn48853 <= z4885_assgn48852;
        z1465_assgn1465 <= z4885_assgn48853;
        z4889_assgn48890 <= z4889_assgn4889;
        z4889_assgn48891 <= z4889_assgn48890;
        z4889_assgn48892 <= z4889_assgn48891;
        z4889_assgn48893 <= z4889_assgn48892;
        z1467_assgn1467 <= z4889_assgn48893;
        z4893_assgn48930 <= z4893_assgn4893;
        z4893_assgn48931 <= z4893_assgn48930;
        z4893_assgn48932 <= z4893_assgn48931;
        z4893_assgn48933 <= z4893_assgn48932;
        z1469_assgn1469 <= z4893_assgn48933;
        z4897_assgn48970 <= z4897_assgn4897;
        z4897_assgn48971 <= z4897_assgn48970;
        z4897_assgn48972 <= z4897_assgn48971;
        z4897_assgn48973 <= z4897_assgn48972;
        z4897_assgn48974 <= z4897_assgn48973;
        z4897_assgn48975 <= z4897_assgn48974;
        z4897_assgn48976 <= z4897_assgn48975;
        z1471_assgn1471 <= z4897_assgn48976;
        z4901_assgn49010 <= z4901_assgn4901;
        z4901_assgn49011 <= z4901_assgn49010;
        z4901_assgn49012 <= z4901_assgn49011;
        z4901_assgn49013 <= z4901_assgn49012;
        z4901_assgn49014 <= z4901_assgn49013;
        z4901_assgn49015 <= z4901_assgn49014;
        z4901_assgn49016 <= z4901_assgn49015;
        z1473_assgn1473 <= z4901_assgn49016;
        z4905_assgn49050 <= z4905_assgn4905;
        z4905_assgn49051 <= z4905_assgn49050;
        z4905_assgn49052 <= z4905_assgn49051;
        z4905_assgn49053 <= z4905_assgn49052;
        z4905_assgn49054 <= z4905_assgn49053;
        z4905_assgn49055 <= z4905_assgn49054;
        z4905_assgn49056 <= z4905_assgn49055;
        z1475_assgn1475 <= z4905_assgn49056;
        z4909_assgn49090 <= z4909_assgn4909;
        z4909_assgn49091 <= z4909_assgn49090;
        z4909_assgn49092 <= z4909_assgn49091;
        z4909_assgn49093 <= z4909_assgn49092;
        z4909_assgn49094 <= z4909_assgn49093;
        z4909_assgn49095 <= z4909_assgn49094;
        z4909_assgn49096 <= z4909_assgn49095;
        z1477_assgn1477 <= z4909_assgn49096;
        z4913_assgn49130 <= z4913_assgn4913;
        z4913_assgn49131 <= z4913_assgn49130;
        z4913_assgn49132 <= z4913_assgn49131;
        z4913_assgn49133 <= z4913_assgn49132;
        z4913_assgn49134 <= z4913_assgn49133;
        z4913_assgn49135 <= z4913_assgn49134;
        z4913_assgn49136 <= z4913_assgn49135;
        z1479_assgn1479 <= z4913_assgn49136;
        z4917_assgn49170 <= z4917_assgn4917;
        z4917_assgn49171 <= z4917_assgn49170;
        z4917_assgn49172 <= z4917_assgn49171;
        z4917_assgn49173 <= z4917_assgn49172;
        z4917_assgn49174 <= z4917_assgn49173;
        z4917_assgn49175 <= z4917_assgn49174;
        z4917_assgn49176 <= z4917_assgn49175;
        z1481_assgn1481 <= z4917_assgn49176;
        z4921_assgn49210 <= z4921_assgn4921;
        z4921_assgn49211 <= z4921_assgn49210;
        z4921_assgn49212 <= z4921_assgn49211;
        z4921_assgn49213 <= z4921_assgn49212;
        z1483_assgn1483 <= z4921_assgn49213;
        z4925_assgn49250 <= z4925_assgn4925;
        z4925_assgn49251 <= z4925_assgn49250;
        z4925_assgn49252 <= z4925_assgn49251;
        z4925_assgn49253 <= z4925_assgn49252;
        z1485_assgn1485 <= z4925_assgn49253;
        z4929_assgn49290 <= z4929_assgn4929;
        z4929_assgn49291 <= z4929_assgn49290;
        z4929_assgn49292 <= z4929_assgn49291;
        z4929_assgn49293 <= z4929_assgn49292;
        z1487_assgn1487 <= z4929_assgn49293;
        z4933_assgn49330 <= z4933_assgn4933;
        z4933_assgn49331 <= z4933_assgn49330;
        z4933_assgn49332 <= z4933_assgn49331;
        z4933_assgn49333 <= z4933_assgn49332;
        z1489_assgn1489 <= z4933_assgn49333;
        z4937_assgn49370 <= z4937_assgn4937;
        z4937_assgn49371 <= z4937_assgn49370;
        z4937_assgn49372 <= z4937_assgn49371;
        z4937_assgn49373 <= z4937_assgn49372;
        z1491_assgn1491 <= z4937_assgn49373;
        z4941_assgn49410 <= z4941_assgn4941;
        z4941_assgn49411 <= z4941_assgn49410;
        z4941_assgn49412 <= z4941_assgn49411;
        z4941_assgn49413 <= z4941_assgn49412;
        z1493_assgn1493 <= z4941_assgn49413;
        c0_G4_mul5_G16_inv0_G256_inv0_reg <= c0_G4_mul5_G16_inv0_G256_inv0;
        d0_G4_mul5_G16_inv0_G256_inv0_reg <= d0_G4_mul5_G16_inv0_G256_inv0;
        c1_G4_mul5_G16_inv0_G256_inv0_reg <= c1_G4_mul5_G16_inv0_G256_inv0;
        d1_G4_mul5_G16_inv0_G256_inv0_reg <= d1_G4_mul5_G16_inv0_G256_inv0;
        z4953_assgn49530 <= z4953_assgn4953;
        z4953_assgn49531 <= z4953_assgn49530;
        z4953_assgn49532 <= z4953_assgn49531;
        z4953_assgn49533 <= z4953_assgn49532;
        z4953_assgn49534 <= z4953_assgn49533;
        z1503_assgn1503 <= z4953_assgn49534;
        z4961_assgn49610 <= z4961_assgn4961;
        z1509_assgn1509 <= z4961_assgn49610;
        z4965_assgn49650 <= z4965_assgn4965;
        z1511_assgn1511 <= z4965_assgn49650;
        cxord_0_G4_mul5_G16_inv0_G256_inv0_reg <= cxord_0_G4_mul5_G16_inv0_G256_inv0;
        r0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
        cxord_1_G4_mul5_G16_inv0_G256_inv0_reg <= cxord_1_G4_mul5_G16_inv0_G256_inv0;
        z4973_assgn49730 <= z4973_assgn4973;
        z1517_assgn1517 <= z4973_assgn49730;
        v1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= v1_hpc20_G4_mul5_G16_inv0_G256_inv0;
        u0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= u0_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p0_hpc20_G4_mul5_G16_inv0_G256_inv0;
        z4983_assgn49830 <= z4983_assgn4983;
        z1525_assgn1525 <= z4983_assgn49830;
        v0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= v0_hpc20_G4_mul5_G16_inv0_G256_inv0;
        u1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= u1_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p3_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p3_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p2_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p2_hpc20_G4_mul5_G16_inv0_G256_inv0;
        z4993_assgn49930 <= z4993_assgn4993;
        z4993_assgn49931 <= z4993_assgn49930;
        z4993_assgn49932 <= z4993_assgn49931;
        z4993_assgn49933 <= z4993_assgn49932;
        z4993_assgn49934 <= z4993_assgn49933;
        z1533_assgn1533 <= z4993_assgn49934;
        z5001_assgn50010 <= z5001_assgn5001;
        z1539_assgn1539 <= z5001_assgn50010;
        z5005_assgn50050 <= z5005_assgn5005;
        z1541_assgn1541 <= z5005_assgn50050;
        z5009_assgn50090 <= z5009_assgn5009;
        z1544_assgn1544 <= z5009_assgn50090;
        r0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
        z5013_assgn50130 <= z5013_assgn5013;
        z1546_assgn1546 <= z5013_assgn50130;
        z5017_assgn50170 <= z5017_assgn5017;
        z5017_assgn50171 <= z5017_assgn50170;
        z1547_assgn1547 <= z5017_assgn50171;
        v1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= v1_hpc21_G4_mul5_G16_inv0_G256_inv0;
        u0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= u0_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p0_hpc21_G4_mul5_G16_inv0_G256_inv0;
        z5027_assgn50270 <= z5027_assgn5027;
        z5027_assgn50271 <= z5027_assgn50270;
        z1555_assgn1555 <= z5027_assgn50271;
        v0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= v0_hpc21_G4_mul5_G16_inv0_G256_inv0;
        u1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= u1_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p3_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p3_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p2_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p2_hpc21_G4_mul5_G16_inv0_G256_inv0;
        z5041_assgn50410 <= z5041_assgn5041;
        z5041_assgn50411 <= z5041_assgn50410;
        z5041_assgn50412 <= z5041_assgn50411;
        z5041_assgn50413 <= z5041_assgn50412;
        z5041_assgn50414 <= z5041_assgn50413;
        z1567_assgn1567 <= z5041_assgn50414;
        z5049_assgn50490 <= z5049_assgn5049;
        z1573_assgn1573 <= z5049_assgn50490;
        z5053_assgn50530 <= z5053_assgn5053;
        z1575_assgn1575 <= z5053_assgn50530;
        z5057_assgn50570 <= z5057_assgn5057;
        z1578_assgn1578 <= z5057_assgn50570;
        r0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
        z5061_assgn50610 <= z5061_assgn5061;
        z1580_assgn1580 <= z5061_assgn50610;
        z5065_assgn50650 <= z5065_assgn5065;
        z5065_assgn50651 <= z5065_assgn50650;
        z1581_assgn1581 <= z5065_assgn50651;
        v1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= v1_hpc22_G4_mul5_G16_inv0_G256_inv0;
        u0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= u0_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p0_hpc22_G4_mul5_G16_inv0_G256_inv0;
        z5075_assgn50750 <= z5075_assgn5075;
        z5075_assgn50751 <= z5075_assgn50750;
        z1589_assgn1589 <= z5075_assgn50751;
        v0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= v0_hpc22_G4_mul5_G16_inv0_G256_inv0;
        u1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= u1_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p3_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p3_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p2_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p2_hpc22_G4_mul5_G16_inv0_G256_inv0;
        z5089_assgn50890 <= z5089_assgn5089;
        z5089_assgn50891 <= z5089_assgn50890;
        z5089_assgn50892 <= z5089_assgn50891;
        z5089_assgn50893 <= z5089_assgn50892;
        z5089_assgn50894 <= z5089_assgn50893;
        z5089_assgn50895 <= z5089_assgn50894;
        z5089_assgn50896 <= z5089_assgn50895;
        z5089_assgn50897 <= z5089_assgn50896;
        z1601_assgn1601 <= z5089_assgn50897;
        z5093_assgn50930 <= z5093_assgn5093;
        z5093_assgn50931 <= z5093_assgn50930;
        z5093_assgn50932 <= z5093_assgn50931;
        z5093_assgn50933 <= z5093_assgn50932;
        z5093_assgn50934 <= z5093_assgn50933;
        z5093_assgn50935 <= z5093_assgn50934;
        z5093_assgn50936 <= z5093_assgn50935;
        z5093_assgn50937 <= z5093_assgn50936;
        z1603_assgn1603 <= z5093_assgn50937;
        z5101_assgn51010 <= z5101_assgn5101;
        z5101_assgn51011 <= z5101_assgn51010;
        z5101_assgn51012 <= z5101_assgn51011;
        z5101_assgn51013 <= z5101_assgn51012;
        z5101_assgn51014 <= z5101_assgn51013;
        z5101_assgn51015 <= z5101_assgn51014;
        z5101_assgn51016 <= z5101_assgn51015;
        z5101_assgn51017 <= z5101_assgn51016;
        z1609_assgn1609 <= z5101_assgn51017;
        z5105_assgn51050 <= z5105_assgn5105;
        z5105_assgn51051 <= z5105_assgn51050;
        z5105_assgn51052 <= z5105_assgn51051;
        z5105_assgn51053 <= z5105_assgn51052;
        z5105_assgn51054 <= z5105_assgn51053;
        z5105_assgn51055 <= z5105_assgn51054;
        z5105_assgn51056 <= z5105_assgn51055;
        z5105_assgn51057 <= z5105_assgn51056;
        z1611_assgn1611 <= z5105_assgn51057;
        z5113_assgn51130 <= z5113_assgn5113;
        z5113_assgn51131 <= z5113_assgn51130;
        z5113_assgn51132 <= z5113_assgn51131;
        z5113_assgn51133 <= z5113_assgn51132;
        z5113_assgn51134 <= z5113_assgn51133;
        z1617_assgn1617 <= z5113_assgn51134;
        z5117_assgn51170 <= z5117_assgn5117;
        z5117_assgn51171 <= z5117_assgn51170;
        z5117_assgn51172 <= z5117_assgn51171;
        z5117_assgn51173 <= z5117_assgn51172;
        z5117_assgn51174 <= z5117_assgn51173;
        z1619_assgn1619 <= z5117_assgn51174;
        z5121_assgn51210 <= z5121_assgn5121;
        z5121_assgn51211 <= z5121_assgn51210;
        z5121_assgn51212 <= z5121_assgn51211;
        z5121_assgn51213 <= z5121_assgn51212;
        z5121_assgn51214 <= z5121_assgn51213;
        z1621_assgn1621 <= z5121_assgn51214;
        z5125_assgn51250 <= z5125_assgn5125;
        z5125_assgn51251 <= z5125_assgn51250;
        z5125_assgn51252 <= z5125_assgn51251;
        z5125_assgn51253 <= z5125_assgn51252;
        z5125_assgn51254 <= z5125_assgn51253;
        z1623_assgn1623 <= z5125_assgn51254;
        z5129_assgn51290 <= z5129_assgn5129;
        z5129_assgn51291 <= z5129_assgn51290;
        z5129_assgn51292 <= z5129_assgn51291;
        z5129_assgn51293 <= z5129_assgn51292;
        z5129_assgn51294 <= z5129_assgn51293;
        z1625_assgn1625 <= z5129_assgn51294;
        z5133_assgn51330 <= z5133_assgn5133;
        z5133_assgn51331 <= z5133_assgn51330;
        z5133_assgn51332 <= z5133_assgn51331;
        z5133_assgn51333 <= z5133_assgn51332;
        z5133_assgn51334 <= z5133_assgn51333;
        z1627_assgn1627 <= z5133_assgn51334;
        z5137_assgn51370 <= z5137_assgn5137;
        z5137_assgn51371 <= z5137_assgn51370;
        z5137_assgn51372 <= z5137_assgn51371;
        z5137_assgn51373 <= z5137_assgn51372;
        z5137_assgn51374 <= z5137_assgn51373;
        z1629_assgn1629 <= z5137_assgn51374;
        z5141_assgn51410 <= z5141_assgn5141;
        z5141_assgn51411 <= z5141_assgn51410;
        z5141_assgn51412 <= z5141_assgn51411;
        z5141_assgn51413 <= z5141_assgn51412;
        z5141_assgn51414 <= z5141_assgn51413;
        z1631_assgn1631 <= z5141_assgn51414;
        z5145_assgn51450 <= z5145_assgn5145;
        z5145_assgn51451 <= z5145_assgn51450;
        z5145_assgn51452 <= z5145_assgn51451;
        z5145_assgn51453 <= z5145_assgn51452;
        z5145_assgn51454 <= z5145_assgn51453;
        z1633_assgn1633 <= z5145_assgn51454;
        z5149_assgn51490 <= z5149_assgn5149;
        z5149_assgn51491 <= z5149_assgn51490;
        z5149_assgn51492 <= z5149_assgn51491;
        z5149_assgn51493 <= z5149_assgn51492;
        z5149_assgn51494 <= z5149_assgn51493;
        z5149_assgn51495 <= z5149_assgn51494;
        z5149_assgn51496 <= z5149_assgn51495;
        z5149_assgn51497 <= z5149_assgn51496;
        z1635_assgn1635 <= z5149_assgn51497;
        z5153_assgn51530 <= z5153_assgn5153;
        z5153_assgn51531 <= z5153_assgn51530;
        z5153_assgn51532 <= z5153_assgn51531;
        z5153_assgn51533 <= z5153_assgn51532;
        z5153_assgn51534 <= z5153_assgn51533;
        z5153_assgn51535 <= z5153_assgn51534;
        z5153_assgn51536 <= z5153_assgn51535;
        z5153_assgn51537 <= z5153_assgn51536;
        z1637_assgn1637 <= z5153_assgn51537;
        z5157_assgn51570 <= z5157_assgn5157;
        z5157_assgn51571 <= z5157_assgn51570;
        z5157_assgn51572 <= z5157_assgn51571;
        z5157_assgn51573 <= z5157_assgn51572;
        z5157_assgn51574 <= z5157_assgn51573;
        z5157_assgn51575 <= z5157_assgn51574;
        z5157_assgn51576 <= z5157_assgn51575;
        z5157_assgn51577 <= z5157_assgn51576;
        z1639_assgn1639 <= z5157_assgn51577;
        z5161_assgn51610 <= z5161_assgn5161;
        z5161_assgn51611 <= z5161_assgn51610;
        z5161_assgn51612 <= z5161_assgn51611;
        z5161_assgn51613 <= z5161_assgn51612;
        z5161_assgn51614 <= z5161_assgn51613;
        z5161_assgn51615 <= z5161_assgn51614;
        z5161_assgn51616 <= z5161_assgn51615;
        z5161_assgn51617 <= z5161_assgn51616;
        z1641_assgn1641 <= z5161_assgn51617;
        z5165_assgn51650 <= z5165_assgn5165;
        z5165_assgn51651 <= z5165_assgn51650;
        z5165_assgn51652 <= z5165_assgn51651;
        z5165_assgn51653 <= z5165_assgn51652;
        z5165_assgn51654 <= z5165_assgn51653;
        z5165_assgn51655 <= z5165_assgn51654;
        z5165_assgn51656 <= z5165_assgn51655;
        z5165_assgn51657 <= z5165_assgn51656;
        z1643_assgn1643 <= z5165_assgn51657;
        z5169_assgn51690 <= z5169_assgn5169;
        z5169_assgn51691 <= z5169_assgn51690;
        z5169_assgn51692 <= z5169_assgn51691;
        z5169_assgn51693 <= z5169_assgn51692;
        z5169_assgn51694 <= z5169_assgn51693;
        z5169_assgn51695 <= z5169_assgn51694;
        z5169_assgn51696 <= z5169_assgn51695;
        z5169_assgn51697 <= z5169_assgn51696;
        z1645_assgn1645 <= z5169_assgn51697;
        z5173_assgn51730 <= z5173_assgn5173;
        z5173_assgn51731 <= z5173_assgn51730;
        z5173_assgn51732 <= z5173_assgn51731;
        z5173_assgn51733 <= z5173_assgn51732;
        z5173_assgn51734 <= z5173_assgn51733;
        z1647_assgn1647 <= z5173_assgn51734;
        z5175_assgn51750 <= z5175_assgn5175;
        z5175_assgn51751 <= z5175_assgn51750;
        z5175_assgn51752 <= z5175_assgn51751;
        z5175_assgn51753 <= z5175_assgn51752;
        z5175_assgn51754 <= z5175_assgn51753;
        z1648_assgn1648 <= z5175_assgn51754;
        z5179_assgn51790 <= z5179_assgn5179;
        z5179_assgn51791 <= z5179_assgn51790;
        z5179_assgn51792 <= z5179_assgn51791;
        z5179_assgn51793 <= z5179_assgn51792;
        z5179_assgn51794 <= z5179_assgn51793;
        z1649_assgn1649 <= z5179_assgn51794;
        z5181_assgn51810 <= z5181_assgn5181;
        z5181_assgn51811 <= z5181_assgn51810;
        z5181_assgn51812 <= z5181_assgn51811;
        z5181_assgn51813 <= z5181_assgn51812;
        z5181_assgn51814 <= z5181_assgn51813;
        z1650_assgn1650 <= z5181_assgn51814;
        z5185_assgn51850 <= z5185_assgn5185;
        z5185_assgn51851 <= z5185_assgn51850;
        z5185_assgn51852 <= z5185_assgn51851;
        z5185_assgn51853 <= z5185_assgn51852;
        z5185_assgn51854 <= z5185_assgn51853;
        z1651_assgn1651 <= z5185_assgn51854;
        z5189_assgn51890 <= z5189_assgn5189;
        z5189_assgn51891 <= z5189_assgn51890;
        z5189_assgn51892 <= z5189_assgn51891;
        z5189_assgn51893 <= z5189_assgn51892;
        z5189_assgn51894 <= z5189_assgn51893;
        z1653_assgn1653 <= z5189_assgn51894;
        z5193_assgn51930 <= z5193_assgn5193;
        z5193_assgn51931 <= z5193_assgn51930;
        z5193_assgn51932 <= z5193_assgn51931;
        z5193_assgn51933 <= z5193_assgn51932;
        z5193_assgn51934 <= z5193_assgn51933;
        z1655_assgn1655 <= z5193_assgn51934;
        z5195_assgn51950 <= z5195_assgn5195;
        z5195_assgn51951 <= z5195_assgn51950;
        z5195_assgn51952 <= z5195_assgn51951;
        z5195_assgn51953 <= z5195_assgn51952;
        z5195_assgn51954 <= z5195_assgn51953;
        z1656_assgn1656 <= z5195_assgn51954;
        z5199_assgn51990 <= z5199_assgn5199;
        z5199_assgn51991 <= z5199_assgn51990;
        z5199_assgn51992 <= z5199_assgn51991;
        z5199_assgn51993 <= z5199_assgn51992;
        z5199_assgn51994 <= z5199_assgn51993;
        z1657_assgn1657 <= z5199_assgn51994;
        z5201_assgn52010 <= z5201_assgn5201;
        z5201_assgn52011 <= z5201_assgn52010;
        z5201_assgn52012 <= z5201_assgn52011;
        z5201_assgn52013 <= z5201_assgn52012;
        z5201_assgn52014 <= z5201_assgn52013;
        z1658_assgn1658 <= z5201_assgn52014;
        z5213_assgn52130 <= z5213_assgn5213;
        z5213_assgn52131 <= z5213_assgn52130;
        z5213_assgn52132 <= z5213_assgn52131;
        z5213_assgn52133 <= z5213_assgn52132;
        z5213_assgn52134 <= z5213_assgn52133;
        z1667_assgn1667 <= z5213_assgn52134;
        z5217_assgn52170 <= z5217_assgn5217;
        z5217_assgn52171 <= z5217_assgn52170;
        z5217_assgn52172 <= z5217_assgn52171;
        z5217_assgn52173 <= z5217_assgn52172;
        z5217_assgn52174 <= z5217_assgn52173;
        z1669_assgn1669 <= z5217_assgn52174;
        z5221_assgn52210 <= z5221_assgn5221;
        z5221_assgn52211 <= z5221_assgn52210;
        z5221_assgn52212 <= z5221_assgn52211;
        z5221_assgn52213 <= z5221_assgn52212;
        z5221_assgn52214 <= z5221_assgn52213;
        z1671_assgn1671 <= z5221_assgn52214;
        z5225_assgn52250 <= z5225_assgn5225;
        z5225_assgn52251 <= z5225_assgn52250;
        z5225_assgn52252 <= z5225_assgn52251;
        z5225_assgn52253 <= z5225_assgn52252;
        z5225_assgn52254 <= z5225_assgn52253;
        z5225_assgn52255 <= z5225_assgn52254;
        z5225_assgn52256 <= z5225_assgn52255;
        z5225_assgn52257 <= z5225_assgn52256;
        z1673_assgn1673 <= z5225_assgn52257;
        z5229_assgn52290 <= z5229_assgn5229;
        z5229_assgn52291 <= z5229_assgn52290;
        z5229_assgn52292 <= z5229_assgn52291;
        z5229_assgn52293 <= z5229_assgn52292;
        z5229_assgn52294 <= z5229_assgn52293;
        z5229_assgn52295 <= z5229_assgn52294;
        z5229_assgn52296 <= z5229_assgn52295;
        z5229_assgn52297 <= z5229_assgn52296;
        z1675_assgn1675 <= z5229_assgn52297;
        z5233_assgn52330 <= z5233_assgn5233;
        z5233_assgn52331 <= z5233_assgn52330;
        z5233_assgn52332 <= z5233_assgn52331;
        z5233_assgn52333 <= z5233_assgn52332;
        z5233_assgn52334 <= z5233_assgn52333;
        z5233_assgn52335 <= z5233_assgn52334;
        z5233_assgn52336 <= z5233_assgn52335;
        z5233_assgn52337 <= z5233_assgn52336;
        z1677_assgn1677 <= z5233_assgn52337;
        z5237_assgn52370 <= z5237_assgn5237;
        z5237_assgn52371 <= z5237_assgn52370;
        z5237_assgn52372 <= z5237_assgn52371;
        z5237_assgn52373 <= z5237_assgn52372;
        z5237_assgn52374 <= z5237_assgn52373;
        z5237_assgn52375 <= z5237_assgn52374;
        z5237_assgn52376 <= z5237_assgn52375;
        z5237_assgn52377 <= z5237_assgn52376;
        z1679_assgn1679 <= z5237_assgn52377;
        z5241_assgn52410 <= z5241_assgn5241;
        z5241_assgn52411 <= z5241_assgn52410;
        z5241_assgn52412 <= z5241_assgn52411;
        z5241_assgn52413 <= z5241_assgn52412;
        z5241_assgn52414 <= z5241_assgn52413;
        z5241_assgn52415 <= z5241_assgn52414;
        z5241_assgn52416 <= z5241_assgn52415;
        z5241_assgn52417 <= z5241_assgn52416;
        z1681_assgn1681 <= z5241_assgn52417;
        z5245_assgn52450 <= z5245_assgn5245;
        z5245_assgn52451 <= z5245_assgn52450;
        z5245_assgn52452 <= z5245_assgn52451;
        z5245_assgn52453 <= z5245_assgn52452;
        z5245_assgn52454 <= z5245_assgn52453;
        z5245_assgn52455 <= z5245_assgn52454;
        z5245_assgn52456 <= z5245_assgn52455;
        z5245_assgn52457 <= z5245_assgn52456;
        z1683_assgn1683 <= z5245_assgn52457;
        z5249_assgn52490 <= z5249_assgn5249;
        z5249_assgn52491 <= z5249_assgn52490;
        z5249_assgn52492 <= z5249_assgn52491;
        z5249_assgn52493 <= z5249_assgn52492;
        z5249_assgn52494 <= z5249_assgn52493;
        z1685_assgn1685 <= z5249_assgn52494;
        z5253_assgn52530 <= z5253_assgn5253;
        z5253_assgn52531 <= z5253_assgn52530;
        z5253_assgn52532 <= z5253_assgn52531;
        z5253_assgn52533 <= z5253_assgn52532;
        z5253_assgn52534 <= z5253_assgn52533;
        z1687_assgn1687 <= z5253_assgn52534;
        z5257_assgn52570 <= z5257_assgn5257;
        z5257_assgn52571 <= z5257_assgn52570;
        z5257_assgn52572 <= z5257_assgn52571;
        z5257_assgn52573 <= z5257_assgn52572;
        z5257_assgn52574 <= z5257_assgn52573;
        z1689_assgn1689 <= z5257_assgn52574;
        z5261_assgn52610 <= z5261_assgn5261;
        z5261_assgn52611 <= z5261_assgn52610;
        z5261_assgn52612 <= z5261_assgn52611;
        z5261_assgn52613 <= z5261_assgn52612;
        z5261_assgn52614 <= z5261_assgn52613;
        z1691_assgn1691 <= z5261_assgn52614;
        z5265_assgn52650 <= z5265_assgn5265;
        z5265_assgn52651 <= z5265_assgn52650;
        z5265_assgn52652 <= z5265_assgn52651;
        z5265_assgn52653 <= z5265_assgn52652;
        z5265_assgn52654 <= z5265_assgn52653;
        z1693_assgn1693 <= z5265_assgn52654;
        z5269_assgn52690 <= z5269_assgn5269;
        z5269_assgn52691 <= z5269_assgn52690;
        z5269_assgn52692 <= z5269_assgn52691;
        z5269_assgn52693 <= z5269_assgn52692;
        z5269_assgn52694 <= z5269_assgn52693;
        z1695_assgn1695 <= z5269_assgn52694;
        c0_G4_mul0_G16_mul1_G256_inv0_reg <= c0_G4_mul0_G16_mul1_G256_inv0;
        d0_G4_mul0_G16_mul1_G256_inv0_reg <= d0_G4_mul0_G16_mul1_G256_inv0;
        c1_G4_mul0_G16_mul1_G256_inv0_reg <= c1_G4_mul0_G16_mul1_G256_inv0;
        d1_G4_mul0_G16_mul1_G256_inv0_reg <= d1_G4_mul0_G16_mul1_G256_inv0;
        z5281_assgn52810 <= z5281_assgn5281;
        z5281_assgn52811 <= z5281_assgn52810;
        z5281_assgn52812 <= z5281_assgn52811;
        z5281_assgn52813 <= z5281_assgn52812;
        z5281_assgn52814 <= z5281_assgn52813;
        z5281_assgn52815 <= z5281_assgn52814;
        z1705_assgn1705 <= z5281_assgn52815;
        z5289_assgn52890 <= z5289_assgn5289;
        z1711_assgn1711 <= z5289_assgn52890;
        z5293_assgn52930 <= z5293_assgn5293;
        z1713_assgn1713 <= z5293_assgn52930;
        cxord_0_G4_mul0_G16_mul1_G256_inv0_reg <= cxord_0_G4_mul0_G16_mul1_G256_inv0;
        r0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
        cxord_1_G4_mul0_G16_mul1_G256_inv0_reg <= cxord_1_G4_mul0_G16_mul1_G256_inv0;
        z5301_assgn53010 <= z5301_assgn5301;
        z1719_assgn1719 <= z5301_assgn53010;
        v1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= v1_hpc20_G4_mul0_G16_mul1_G256_inv0;
        u0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= u0_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p0_hpc20_G4_mul0_G16_mul1_G256_inv0;
        z5311_assgn53110 <= z5311_assgn5311;
        z1727_assgn1727 <= z5311_assgn53110;
        v0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= v0_hpc20_G4_mul0_G16_mul1_G256_inv0;
        u1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= u1_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p3_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p3_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p2_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p2_hpc20_G4_mul0_G16_mul1_G256_inv0;
        z5321_assgn53210 <= z5321_assgn5321;
        z5321_assgn53211 <= z5321_assgn53210;
        z5321_assgn53212 <= z5321_assgn53211;
        z5321_assgn53213 <= z5321_assgn53212;
        z5321_assgn53214 <= z5321_assgn53213;
        z5321_assgn53215 <= z5321_assgn53214;
        z1735_assgn1735 <= z5321_assgn53215;
        z5329_assgn53290 <= z5329_assgn5329;
        z1741_assgn1741 <= z5329_assgn53290;
        z5333_assgn53330 <= z5333_assgn5333;
        z1743_assgn1743 <= z5333_assgn53330;
        z5337_assgn53370 <= z5337_assgn5337;
        z1746_assgn1746 <= z5337_assgn53370;
        r0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
        z5341_assgn53410 <= z5341_assgn5341;
        z1748_assgn1748 <= z5341_assgn53410;
        z5345_assgn53450 <= z5345_assgn5345;
        z5345_assgn53451 <= z5345_assgn53450;
        z1749_assgn1749 <= z5345_assgn53451;
        v1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= v1_hpc21_G4_mul0_G16_mul1_G256_inv0;
        u0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= u0_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p0_hpc21_G4_mul0_G16_mul1_G256_inv0;
        z5355_assgn53550 <= z5355_assgn5355;
        z5355_assgn53551 <= z5355_assgn53550;
        z1757_assgn1757 <= z5355_assgn53551;
        v0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= v0_hpc21_G4_mul0_G16_mul1_G256_inv0;
        u1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= u1_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p3_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p3_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p2_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p2_hpc21_G4_mul0_G16_mul1_G256_inv0;
        z5369_assgn53690 <= z5369_assgn5369;
        z5369_assgn53691 <= z5369_assgn53690;
        z5369_assgn53692 <= z5369_assgn53691;
        z5369_assgn53693 <= z5369_assgn53692;
        z5369_assgn53694 <= z5369_assgn53693;
        z5369_assgn53695 <= z5369_assgn53694;
        z1769_assgn1769 <= z5369_assgn53695;
        z5377_assgn53770 <= z5377_assgn5377;
        z1775_assgn1775 <= z5377_assgn53770;
        z5381_assgn53810 <= z5381_assgn5381;
        z1777_assgn1777 <= z5381_assgn53810;
        z5385_assgn53850 <= z5385_assgn5385;
        z1780_assgn1780 <= z5385_assgn53850;
        r0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
        z5389_assgn53890 <= z5389_assgn5389;
        z1782_assgn1782 <= z5389_assgn53890;
        z5393_assgn53930 <= z5393_assgn5393;
        z5393_assgn53931 <= z5393_assgn53930;
        z1783_assgn1783 <= z5393_assgn53931;
        v1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= v1_hpc22_G4_mul0_G16_mul1_G256_inv0;
        u0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= u0_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p0_hpc22_G4_mul0_G16_mul1_G256_inv0;
        z5403_assgn54030 <= z5403_assgn5403;
        z5403_assgn54031 <= z5403_assgn54030;
        z1791_assgn1791 <= z5403_assgn54031;
        v0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= v0_hpc22_G4_mul0_G16_mul1_G256_inv0;
        u1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= u1_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p3_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p3_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p2_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p2_hpc22_G4_mul0_G16_mul1_G256_inv0;
        z5417_assgn54170 <= z5417_assgn5417;
        z5417_assgn54171 <= z5417_assgn54170;
        z5417_assgn54172 <= z5417_assgn54171;
        z5417_assgn54173 <= z5417_assgn54172;
        z5417_assgn54174 <= z5417_assgn54173;
        z5417_assgn54175 <= z5417_assgn54174;
        z5417_assgn54176 <= z5417_assgn54175;
        z5417_assgn54177 <= z5417_assgn54176;
        z5417_assgn54178 <= z5417_assgn54177;
        z1803_assgn1803 <= z5417_assgn54178;
        z5421_assgn54210 <= z5421_assgn5421;
        z5421_assgn54211 <= z5421_assgn54210;
        z5421_assgn54212 <= z5421_assgn54211;
        z5421_assgn54213 <= z5421_assgn54212;
        z5421_assgn54214 <= z5421_assgn54213;
        z5421_assgn54215 <= z5421_assgn54214;
        z5421_assgn54216 <= z5421_assgn54215;
        z5421_assgn54217 <= z5421_assgn54216;
        z5421_assgn54218 <= z5421_assgn54217;
        z1805_assgn1805 <= z5421_assgn54218;
        z5429_assgn54290 <= z5429_assgn5429;
        z5429_assgn54291 <= z5429_assgn54290;
        z5429_assgn54292 <= z5429_assgn54291;
        z5429_assgn54293 <= z5429_assgn54292;
        z5429_assgn54294 <= z5429_assgn54293;
        z5429_assgn54295 <= z5429_assgn54294;
        z5429_assgn54296 <= z5429_assgn54295;
        z5429_assgn54297 <= z5429_assgn54296;
        z5429_assgn54298 <= z5429_assgn54297;
        z1811_assgn1811 <= z5429_assgn54298;
        z5433_assgn54330 <= z5433_assgn5433;
        z5433_assgn54331 <= z5433_assgn54330;
        z5433_assgn54332 <= z5433_assgn54331;
        z5433_assgn54333 <= z5433_assgn54332;
        z5433_assgn54334 <= z5433_assgn54333;
        z5433_assgn54335 <= z5433_assgn54334;
        z5433_assgn54336 <= z5433_assgn54335;
        z5433_assgn54337 <= z5433_assgn54336;
        z5433_assgn54338 <= z5433_assgn54337;
        z1813_assgn1813 <= z5433_assgn54338;
        z5437_assgn54370 <= z5437_assgn5437;
        z5437_assgn54371 <= z5437_assgn54370;
        z5437_assgn54372 <= z5437_assgn54371;
        z5437_assgn54373 <= z5437_assgn54372;
        z5437_assgn54374 <= z5437_assgn54373;
        z5437_assgn54375 <= z5437_assgn54374;
        z5437_assgn54376 <= z5437_assgn54375;
        z5437_assgn54377 <= z5437_assgn54376;
        z5437_assgn54378 <= z5437_assgn54377;
        z1815_assgn1815 <= z5437_assgn54378;
        z5441_assgn54410 <= z5441_assgn5441;
        z5441_assgn54411 <= z5441_assgn54410;
        z5441_assgn54412 <= z5441_assgn54411;
        z5441_assgn54413 <= z5441_assgn54412;
        z5441_assgn54414 <= z5441_assgn54413;
        z5441_assgn54415 <= z5441_assgn54414;
        z5441_assgn54416 <= z5441_assgn54415;
        z5441_assgn54417 <= z5441_assgn54416;
        z5441_assgn54418 <= z5441_assgn54417;
        z1817_assgn1817 <= z5441_assgn54418;
        z5445_assgn54450 <= z5445_assgn5445;
        z5445_assgn54451 <= z5445_assgn54450;
        z5445_assgn54452 <= z5445_assgn54451;
        z5445_assgn54453 <= z5445_assgn54452;
        z5445_assgn54454 <= z5445_assgn54453;
        z5445_assgn54455 <= z5445_assgn54454;
        z5445_assgn54456 <= z5445_assgn54455;
        z5445_assgn54457 <= z5445_assgn54456;
        z5445_assgn54458 <= z5445_assgn54457;
        z1819_assgn1819 <= z5445_assgn54458;
        z5449_assgn54490 <= z5449_assgn5449;
        z5449_assgn54491 <= z5449_assgn54490;
        z5449_assgn54492 <= z5449_assgn54491;
        z5449_assgn54493 <= z5449_assgn54492;
        z5449_assgn54494 <= z5449_assgn54493;
        z5449_assgn54495 <= z5449_assgn54494;
        z5449_assgn54496 <= z5449_assgn54495;
        z5449_assgn54497 <= z5449_assgn54496;
        z5449_assgn54498 <= z5449_assgn54497;
        z1821_assgn1821 <= z5449_assgn54498;
        z5461_assgn54610 <= z5461_assgn5461;
        z5461_assgn54611 <= z5461_assgn54610;
        z5461_assgn54612 <= z5461_assgn54611;
        z5461_assgn54613 <= z5461_assgn54612;
        z5461_assgn54614 <= z5461_assgn54613;
        z5461_assgn54615 <= z5461_assgn54614;
        z5461_assgn54616 <= z5461_assgn54615;
        z5461_assgn54617 <= z5461_assgn54616;
        z5461_assgn54618 <= z5461_assgn54617;
        z1831_assgn1831 <= z5461_assgn54618;
        z5465_assgn54650 <= z5465_assgn5465;
        z5465_assgn54651 <= z5465_assgn54650;
        z5465_assgn54652 <= z5465_assgn54651;
        z5465_assgn54653 <= z5465_assgn54652;
        z5465_assgn54654 <= z5465_assgn54653;
        z5465_assgn54655 <= z5465_assgn54654;
        z5465_assgn54656 <= z5465_assgn54655;
        z5465_assgn54657 <= z5465_assgn54656;
        z5465_assgn54658 <= z5465_assgn54657;
        z1833_assgn1833 <= z5465_assgn54658;
        z5473_assgn54730 <= z5473_assgn5473;
        z5473_assgn54731 <= z5473_assgn54730;
        z5473_assgn54732 <= z5473_assgn54731;
        z5473_assgn54733 <= z5473_assgn54732;
        z5473_assgn54734 <= z5473_assgn54733;
        z1839_assgn1839 <= z5473_assgn54734;
        z5477_assgn54770 <= z5477_assgn5477;
        z5477_assgn54771 <= z5477_assgn54770;
        z5477_assgn54772 <= z5477_assgn54771;
        z5477_assgn54773 <= z5477_assgn54772;
        z5477_assgn54774 <= z5477_assgn54773;
        z1841_assgn1841 <= z5477_assgn54774;
        z5481_assgn54810 <= z5481_assgn5481;
        z5481_assgn54811 <= z5481_assgn54810;
        z5481_assgn54812 <= z5481_assgn54811;
        z5481_assgn54813 <= z5481_assgn54812;
        z5481_assgn54814 <= z5481_assgn54813;
        z1843_assgn1843 <= z5481_assgn54814;
        z5485_assgn54850 <= z5485_assgn5485;
        z5485_assgn54851 <= z5485_assgn54850;
        z5485_assgn54852 <= z5485_assgn54851;
        z5485_assgn54853 <= z5485_assgn54852;
        z5485_assgn54854 <= z5485_assgn54853;
        z5485_assgn54855 <= z5485_assgn54854;
        z5485_assgn54856 <= z5485_assgn54855;
        z5485_assgn54857 <= z5485_assgn54856;
        z1845_assgn1845 <= z5485_assgn54857;
        z5489_assgn54890 <= z5489_assgn5489;
        z5489_assgn54891 <= z5489_assgn54890;
        z5489_assgn54892 <= z5489_assgn54891;
        z5489_assgn54893 <= z5489_assgn54892;
        z5489_assgn54894 <= z5489_assgn54893;
        z5489_assgn54895 <= z5489_assgn54894;
        z5489_assgn54896 <= z5489_assgn54895;
        z5489_assgn54897 <= z5489_assgn54896;
        z1847_assgn1847 <= z5489_assgn54897;
        z5493_assgn54930 <= z5493_assgn5493;
        z5493_assgn54931 <= z5493_assgn54930;
        z5493_assgn54932 <= z5493_assgn54931;
        z5493_assgn54933 <= z5493_assgn54932;
        z5493_assgn54934 <= z5493_assgn54933;
        z5493_assgn54935 <= z5493_assgn54934;
        z5493_assgn54936 <= z5493_assgn54935;
        z5493_assgn54937 <= z5493_assgn54936;
        z1849_assgn1849 <= z5493_assgn54937;
        z5497_assgn54970 <= z5497_assgn5497;
        z5497_assgn54971 <= z5497_assgn54970;
        z5497_assgn54972 <= z5497_assgn54971;
        z5497_assgn54973 <= z5497_assgn54972;
        z5497_assgn54974 <= z5497_assgn54973;
        z5497_assgn54975 <= z5497_assgn54974;
        z5497_assgn54976 <= z5497_assgn54975;
        z5497_assgn54977 <= z5497_assgn54976;
        z1851_assgn1851 <= z5497_assgn54977;
        z5501_assgn55010 <= z5501_assgn5501;
        z5501_assgn55011 <= z5501_assgn55010;
        z5501_assgn55012 <= z5501_assgn55011;
        z5501_assgn55013 <= z5501_assgn55012;
        z5501_assgn55014 <= z5501_assgn55013;
        z5501_assgn55015 <= z5501_assgn55014;
        z5501_assgn55016 <= z5501_assgn55015;
        z5501_assgn55017 <= z5501_assgn55016;
        z1853_assgn1853 <= z5501_assgn55017;
        z5505_assgn55050 <= z5505_assgn5505;
        z5505_assgn55051 <= z5505_assgn55050;
        z5505_assgn55052 <= z5505_assgn55051;
        z5505_assgn55053 <= z5505_assgn55052;
        z5505_assgn55054 <= z5505_assgn55053;
        z5505_assgn55055 <= z5505_assgn55054;
        z5505_assgn55056 <= z5505_assgn55055;
        z5505_assgn55057 <= z5505_assgn55056;
        z1855_assgn1855 <= z5505_assgn55057;
        z5509_assgn55090 <= z5509_assgn5509;
        z5509_assgn55091 <= z5509_assgn55090;
        z5509_assgn55092 <= z5509_assgn55091;
        z5509_assgn55093 <= z5509_assgn55092;
        z5509_assgn55094 <= z5509_assgn55093;
        z1857_assgn1857 <= z5509_assgn55094;
        z5513_assgn55130 <= z5513_assgn5513;
        z5513_assgn55131 <= z5513_assgn55130;
        z5513_assgn55132 <= z5513_assgn55131;
        z5513_assgn55133 <= z5513_assgn55132;
        z5513_assgn55134 <= z5513_assgn55133;
        z1859_assgn1859 <= z5513_assgn55134;
        z5517_assgn55170 <= z5517_assgn5517;
        z5517_assgn55171 <= z5517_assgn55170;
        z5517_assgn55172 <= z5517_assgn55171;
        z5517_assgn55173 <= z5517_assgn55172;
        z5517_assgn55174 <= z5517_assgn55173;
        z1861_assgn1861 <= z5517_assgn55174;
        z5521_assgn55210 <= z5521_assgn5521;
        z5521_assgn55211 <= z5521_assgn55210;
        z5521_assgn55212 <= z5521_assgn55211;
        z5521_assgn55213 <= z5521_assgn55212;
        z5521_assgn55214 <= z5521_assgn55213;
        z1863_assgn1863 <= z5521_assgn55214;
        z5525_assgn55250 <= z5525_assgn5525;
        z5525_assgn55251 <= z5525_assgn55250;
        z5525_assgn55252 <= z5525_assgn55251;
        z5525_assgn55253 <= z5525_assgn55252;
        z5525_assgn55254 <= z5525_assgn55253;
        z1865_assgn1865 <= z5525_assgn55254;
        z5529_assgn55290 <= z5529_assgn5529;
        z5529_assgn55291 <= z5529_assgn55290;
        z5529_assgn55292 <= z5529_assgn55291;
        z5529_assgn55293 <= z5529_assgn55292;
        z5529_assgn55294 <= z5529_assgn55293;
        z1867_assgn1867 <= z5529_assgn55294;
        c0_G4_mul1_G16_mul1_G256_inv0_reg <= c0_G4_mul1_G16_mul1_G256_inv0;
        d0_G4_mul1_G16_mul1_G256_inv0_reg <= d0_G4_mul1_G16_mul1_G256_inv0;
        c1_G4_mul1_G16_mul1_G256_inv0_reg <= c1_G4_mul1_G16_mul1_G256_inv0;
        d1_G4_mul1_G16_mul1_G256_inv0_reg <= d1_G4_mul1_G16_mul1_G256_inv0;
        z5541_assgn55410 <= z5541_assgn5541;
        z5541_assgn55411 <= z5541_assgn55410;
        z5541_assgn55412 <= z5541_assgn55411;
        z5541_assgn55413 <= z5541_assgn55412;
        z5541_assgn55414 <= z5541_assgn55413;
        z5541_assgn55415 <= z5541_assgn55414;
        z1877_assgn1877 <= z5541_assgn55415;
        z5549_assgn55490 <= z5549_assgn5549;
        z1883_assgn1883 <= z5549_assgn55490;
        z5553_assgn55530 <= z5553_assgn5553;
        z1885_assgn1885 <= z5553_assgn55530;
        cxord_0_G4_mul1_G16_mul1_G256_inv0_reg <= cxord_0_G4_mul1_G16_mul1_G256_inv0;
        r0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
        cxord_1_G4_mul1_G16_mul1_G256_inv0_reg <= cxord_1_G4_mul1_G16_mul1_G256_inv0;
        z5561_assgn55610 <= z5561_assgn5561;
        z1891_assgn1891 <= z5561_assgn55610;
        v1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= v1_hpc20_G4_mul1_G16_mul1_G256_inv0;
        u0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= u0_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p0_hpc20_G4_mul1_G16_mul1_G256_inv0;
        z5571_assgn55710 <= z5571_assgn5571;
        z1899_assgn1899 <= z5571_assgn55710;
        v0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= v0_hpc20_G4_mul1_G16_mul1_G256_inv0;
        u1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= u1_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p3_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p3_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p2_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p2_hpc20_G4_mul1_G16_mul1_G256_inv0;
        z5581_assgn55810 <= z5581_assgn5581;
        z5581_assgn55811 <= z5581_assgn55810;
        z5581_assgn55812 <= z5581_assgn55811;
        z5581_assgn55813 <= z5581_assgn55812;
        z5581_assgn55814 <= z5581_assgn55813;
        z5581_assgn55815 <= z5581_assgn55814;
        z1907_assgn1907 <= z5581_assgn55815;
        z5589_assgn55890 <= z5589_assgn5589;
        z1913_assgn1913 <= z5589_assgn55890;
        z5593_assgn55930 <= z5593_assgn5593;
        z1915_assgn1915 <= z5593_assgn55930;
        z5597_assgn55970 <= z5597_assgn5597;
        z1918_assgn1918 <= z5597_assgn55970;
        r0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
        z5601_assgn56010 <= z5601_assgn5601;
        z1920_assgn1920 <= z5601_assgn56010;
        z5605_assgn56050 <= z5605_assgn5605;
        z5605_assgn56051 <= z5605_assgn56050;
        z1921_assgn1921 <= z5605_assgn56051;
        v1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= v1_hpc21_G4_mul1_G16_mul1_G256_inv0;
        u0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= u0_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p0_hpc21_G4_mul1_G16_mul1_G256_inv0;
        z5615_assgn56150 <= z5615_assgn5615;
        z5615_assgn56151 <= z5615_assgn56150;
        z1929_assgn1929 <= z5615_assgn56151;
        v0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= v0_hpc21_G4_mul1_G16_mul1_G256_inv0;
        u1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= u1_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p3_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p3_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p2_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p2_hpc21_G4_mul1_G16_mul1_G256_inv0;
        z5629_assgn56290 <= z5629_assgn5629;
        z5629_assgn56291 <= z5629_assgn56290;
        z5629_assgn56292 <= z5629_assgn56291;
        z5629_assgn56293 <= z5629_assgn56292;
        z5629_assgn56294 <= z5629_assgn56293;
        z5629_assgn56295 <= z5629_assgn56294;
        z1941_assgn1941 <= z5629_assgn56295;
        z5637_assgn56370 <= z5637_assgn5637;
        z1947_assgn1947 <= z5637_assgn56370;
        z5641_assgn56410 <= z5641_assgn5641;
        z1949_assgn1949 <= z5641_assgn56410;
        z5645_assgn56450 <= z5645_assgn5645;
        z1952_assgn1952 <= z5645_assgn56450;
        r0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
        z5649_assgn56490 <= z5649_assgn5649;
        z1954_assgn1954 <= z5649_assgn56490;
        z5653_assgn56530 <= z5653_assgn5653;
        z5653_assgn56531 <= z5653_assgn56530;
        z1955_assgn1955 <= z5653_assgn56531;
        v1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= v1_hpc22_G4_mul1_G16_mul1_G256_inv0;
        u0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= u0_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p0_hpc22_G4_mul1_G16_mul1_G256_inv0;
        z5663_assgn56630 <= z5663_assgn5663;
        z5663_assgn56631 <= z5663_assgn56630;
        z1963_assgn1963 <= z5663_assgn56631;
        v0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= v0_hpc22_G4_mul1_G16_mul1_G256_inv0;
        u1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= u1_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p3_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p3_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p2_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p2_hpc22_G4_mul1_G16_mul1_G256_inv0;
        z5677_assgn56770 <= z5677_assgn5677;
        z5677_assgn56771 <= z5677_assgn56770;
        z5677_assgn56772 <= z5677_assgn56771;
        z5677_assgn56773 <= z5677_assgn56772;
        z5677_assgn56774 <= z5677_assgn56773;
        z5677_assgn56775 <= z5677_assgn56774;
        z5677_assgn56776 <= z5677_assgn56775;
        z5677_assgn56777 <= z5677_assgn56776;
        z5677_assgn56778 <= z5677_assgn56777;
        z1975_assgn1975 <= z5677_assgn56778;
        z5681_assgn56810 <= z5681_assgn5681;
        z5681_assgn56811 <= z5681_assgn56810;
        z5681_assgn56812 <= z5681_assgn56811;
        z5681_assgn56813 <= z5681_assgn56812;
        z5681_assgn56814 <= z5681_assgn56813;
        z5681_assgn56815 <= z5681_assgn56814;
        z5681_assgn56816 <= z5681_assgn56815;
        z5681_assgn56817 <= z5681_assgn56816;
        z5681_assgn56818 <= z5681_assgn56817;
        z1977_assgn1977 <= z5681_assgn56818;
        z5693_assgn56930 <= z5693_assgn5693;
        z5693_assgn56931 <= z5693_assgn56930;
        z5693_assgn56932 <= z5693_assgn56931;
        z5693_assgn56933 <= z5693_assgn56932;
        z5693_assgn56934 <= z5693_assgn56933;
        z1987_assgn1987 <= z5693_assgn56934;
        z5697_assgn56970 <= z5697_assgn5697;
        z5697_assgn56971 <= z5697_assgn56970;
        z5697_assgn56972 <= z5697_assgn56971;
        z5697_assgn56973 <= z5697_assgn56972;
        z5697_assgn56974 <= z5697_assgn56973;
        z1989_assgn1989 <= z5697_assgn56974;
        z5701_assgn57010 <= z5701_assgn5701;
        z5701_assgn57011 <= z5701_assgn57010;
        z5701_assgn57012 <= z5701_assgn57011;
        z5701_assgn57013 <= z5701_assgn57012;
        z5701_assgn57014 <= z5701_assgn57013;
        z1991_assgn1991 <= z5701_assgn57014;
        z5705_assgn57050 <= z5705_assgn5705;
        z5705_assgn57051 <= z5705_assgn57050;
        z5705_assgn57052 <= z5705_assgn57051;
        z5705_assgn57053 <= z5705_assgn57052;
        z5705_assgn57054 <= z5705_assgn57053;
        z5705_assgn57055 <= z5705_assgn57054;
        z5705_assgn57056 <= z5705_assgn57055;
        z5705_assgn57057 <= z5705_assgn57056;
        z1993_assgn1993 <= z5705_assgn57057;
        z5709_assgn57090 <= z5709_assgn5709;
        z5709_assgn57091 <= z5709_assgn57090;
        z5709_assgn57092 <= z5709_assgn57091;
        z5709_assgn57093 <= z5709_assgn57092;
        z5709_assgn57094 <= z5709_assgn57093;
        z5709_assgn57095 <= z5709_assgn57094;
        z5709_assgn57096 <= z5709_assgn57095;
        z5709_assgn57097 <= z5709_assgn57096;
        z1995_assgn1995 <= z5709_assgn57097;
        z5713_assgn57130 <= z5713_assgn5713;
        z5713_assgn57131 <= z5713_assgn57130;
        z5713_assgn57132 <= z5713_assgn57131;
        z5713_assgn57133 <= z5713_assgn57132;
        z5713_assgn57134 <= z5713_assgn57133;
        z5713_assgn57135 <= z5713_assgn57134;
        z5713_assgn57136 <= z5713_assgn57135;
        z5713_assgn57137 <= z5713_assgn57136;
        z1997_assgn1997 <= z5713_assgn57137;
        z5717_assgn57170 <= z5717_assgn5717;
        z5717_assgn57171 <= z5717_assgn57170;
        z5717_assgn57172 <= z5717_assgn57171;
        z5717_assgn57173 <= z5717_assgn57172;
        z5717_assgn57174 <= z5717_assgn57173;
        z5717_assgn57175 <= z5717_assgn57174;
        z5717_assgn57176 <= z5717_assgn57175;
        z5717_assgn57177 <= z5717_assgn57176;
        z1999_assgn1999 <= z5717_assgn57177;
        z5721_assgn57210 <= z5721_assgn5721;
        z5721_assgn57211 <= z5721_assgn57210;
        z5721_assgn57212 <= z5721_assgn57211;
        z5721_assgn57213 <= z5721_assgn57212;
        z5721_assgn57214 <= z5721_assgn57213;
        z5721_assgn57215 <= z5721_assgn57214;
        z5721_assgn57216 <= z5721_assgn57215;
        z5721_assgn57217 <= z5721_assgn57216;
        z2001_assgn2001 <= z5721_assgn57217;
        z5725_assgn57250 <= z5725_assgn5725;
        z5725_assgn57251 <= z5725_assgn57250;
        z5725_assgn57252 <= z5725_assgn57251;
        z5725_assgn57253 <= z5725_assgn57252;
        z5725_assgn57254 <= z5725_assgn57253;
        z5725_assgn57255 <= z5725_assgn57254;
        z5725_assgn57256 <= z5725_assgn57255;
        z5725_assgn57257 <= z5725_assgn57256;
        z2003_assgn2003 <= z5725_assgn57257;
        z5729_assgn57290 <= z5729_assgn5729;
        z5729_assgn57291 <= z5729_assgn57290;
        z5729_assgn57292 <= z5729_assgn57291;
        z5729_assgn57293 <= z5729_assgn57292;
        z5729_assgn57294 <= z5729_assgn57293;
        z2005_assgn2005 <= z5729_assgn57294;
        z5733_assgn57330 <= z5733_assgn5733;
        z5733_assgn57331 <= z5733_assgn57330;
        z5733_assgn57332 <= z5733_assgn57331;
        z5733_assgn57333 <= z5733_assgn57332;
        z5733_assgn57334 <= z5733_assgn57333;
        z2007_assgn2007 <= z5733_assgn57334;
        z5737_assgn57370 <= z5737_assgn5737;
        z5737_assgn57371 <= z5737_assgn57370;
        z5737_assgn57372 <= z5737_assgn57371;
        z5737_assgn57373 <= z5737_assgn57372;
        z5737_assgn57374 <= z5737_assgn57373;
        z2009_assgn2009 <= z5737_assgn57374;
        z5741_assgn57410 <= z5741_assgn5741;
        z5741_assgn57411 <= z5741_assgn57410;
        z5741_assgn57412 <= z5741_assgn57411;
        z5741_assgn57413 <= z5741_assgn57412;
        z5741_assgn57414 <= z5741_assgn57413;
        z2011_assgn2011 <= z5741_assgn57414;
        z5745_assgn57450 <= z5745_assgn5745;
        z5745_assgn57451 <= z5745_assgn57450;
        z5745_assgn57452 <= z5745_assgn57451;
        z5745_assgn57453 <= z5745_assgn57452;
        z5745_assgn57454 <= z5745_assgn57453;
        z2013_assgn2013 <= z5745_assgn57454;
        z5749_assgn57490 <= z5749_assgn5749;
        z5749_assgn57491 <= z5749_assgn57490;
        z5749_assgn57492 <= z5749_assgn57491;
        z5749_assgn57493 <= z5749_assgn57492;
        z5749_assgn57494 <= z5749_assgn57493;
        z2015_assgn2015 <= z5749_assgn57494;
        c0_G4_mul2_G16_mul1_G256_inv0_reg <= c0_G4_mul2_G16_mul1_G256_inv0;
        d0_G4_mul2_G16_mul1_G256_inv0_reg <= d0_G4_mul2_G16_mul1_G256_inv0;
        c1_G4_mul2_G16_mul1_G256_inv0_reg <= c1_G4_mul2_G16_mul1_G256_inv0;
        d1_G4_mul2_G16_mul1_G256_inv0_reg <= d1_G4_mul2_G16_mul1_G256_inv0;
        z5761_assgn57610 <= z5761_assgn5761;
        z5761_assgn57611 <= z5761_assgn57610;
        z5761_assgn57612 <= z5761_assgn57611;
        z5761_assgn57613 <= z5761_assgn57612;
        z5761_assgn57614 <= z5761_assgn57613;
        z5761_assgn57615 <= z5761_assgn57614;
        z2025_assgn2025 <= z5761_assgn57615;
        z5769_assgn57690 <= z5769_assgn5769;
        z2031_assgn2031 <= z5769_assgn57690;
        z5773_assgn57730 <= z5773_assgn5773;
        z2033_assgn2033 <= z5773_assgn57730;
        cxord_0_G4_mul2_G16_mul1_G256_inv0_reg <= cxord_0_G4_mul2_G16_mul1_G256_inv0;
        r0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
        cxord_1_G4_mul2_G16_mul1_G256_inv0_reg <= cxord_1_G4_mul2_G16_mul1_G256_inv0;
        z5781_assgn57810 <= z5781_assgn5781;
        z2039_assgn2039 <= z5781_assgn57810;
        v1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= v1_hpc20_G4_mul2_G16_mul1_G256_inv0;
        u0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= u0_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p0_hpc20_G4_mul2_G16_mul1_G256_inv0;
        z5791_assgn57910 <= z5791_assgn5791;
        z2047_assgn2047 <= z5791_assgn57910;
        v0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= v0_hpc20_G4_mul2_G16_mul1_G256_inv0;
        u1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= u1_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p3_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p3_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p2_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p2_hpc20_G4_mul2_G16_mul1_G256_inv0;
        z5801_assgn58010 <= z5801_assgn5801;
        z5801_assgn58011 <= z5801_assgn58010;
        z5801_assgn58012 <= z5801_assgn58011;
        z5801_assgn58013 <= z5801_assgn58012;
        z5801_assgn58014 <= z5801_assgn58013;
        z5801_assgn58015 <= z5801_assgn58014;
        z2055_assgn2055 <= z5801_assgn58015;
        z5809_assgn58090 <= z5809_assgn5809;
        z2061_assgn2061 <= z5809_assgn58090;
        z5813_assgn58130 <= z5813_assgn5813;
        z2063_assgn2063 <= z5813_assgn58130;
        z5817_assgn58170 <= z5817_assgn5817;
        z2066_assgn2066 <= z5817_assgn58170;
        r0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
        z5821_assgn58210 <= z5821_assgn5821;
        z2068_assgn2068 <= z5821_assgn58210;
        z5825_assgn58250 <= z5825_assgn5825;
        z5825_assgn58251 <= z5825_assgn58250;
        z2069_assgn2069 <= z5825_assgn58251;
        v1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= v1_hpc21_G4_mul2_G16_mul1_G256_inv0;
        u0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= u0_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p0_hpc21_G4_mul2_G16_mul1_G256_inv0;
        z5835_assgn58350 <= z5835_assgn5835;
        z5835_assgn58351 <= z5835_assgn58350;
        z2077_assgn2077 <= z5835_assgn58351;
        v0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= v0_hpc21_G4_mul2_G16_mul1_G256_inv0;
        u1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= u1_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p3_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p3_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p2_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p2_hpc21_G4_mul2_G16_mul1_G256_inv0;
        z5849_assgn58490 <= z5849_assgn5849;
        z5849_assgn58491 <= z5849_assgn58490;
        z5849_assgn58492 <= z5849_assgn58491;
        z5849_assgn58493 <= z5849_assgn58492;
        z5849_assgn58494 <= z5849_assgn58493;
        z5849_assgn58495 <= z5849_assgn58494;
        z2089_assgn2089 <= z5849_assgn58495;
        z5857_assgn58570 <= z5857_assgn5857;
        z2095_assgn2095 <= z5857_assgn58570;
        z5861_assgn58610 <= z5861_assgn5861;
        z2097_assgn2097 <= z5861_assgn58610;
        z5865_assgn58650 <= z5865_assgn5865;
        z2100_assgn2100 <= z5865_assgn58650;
        r0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
        z5869_assgn58690 <= z5869_assgn5869;
        z2102_assgn2102 <= z5869_assgn58690;
        z5873_assgn58730 <= z5873_assgn5873;
        z5873_assgn58731 <= z5873_assgn58730;
        z2103_assgn2103 <= z5873_assgn58731;
        v1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= v1_hpc22_G4_mul2_G16_mul1_G256_inv0;
        u0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= u0_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p0_hpc22_G4_mul2_G16_mul1_G256_inv0;
        z5883_assgn58830 <= z5883_assgn5883;
        z5883_assgn58831 <= z5883_assgn58830;
        z2111_assgn2111 <= z5883_assgn58831;
        v0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= v0_hpc22_G4_mul2_G16_mul1_G256_inv0;
        u1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= u1_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p3_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p3_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p2_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p2_hpc22_G4_mul2_G16_mul1_G256_inv0;
        z5897_assgn58970 <= z5897_assgn5897;
        z5897_assgn58971 <= z5897_assgn58970;
        z5897_assgn58972 <= z5897_assgn58971;
        z5897_assgn58973 <= z5897_assgn58972;
        z5897_assgn58974 <= z5897_assgn58973;
        z5897_assgn58975 <= z5897_assgn58974;
        z5897_assgn58976 <= z5897_assgn58975;
        z5897_assgn58977 <= z5897_assgn58976;
        z5897_assgn58978 <= z5897_assgn58977;
        z2123_assgn2123 <= z5897_assgn58978;
        z5901_assgn59010 <= z5901_assgn5901;
        z5901_assgn59011 <= z5901_assgn59010;
        z5901_assgn59012 <= z5901_assgn59011;
        z5901_assgn59013 <= z5901_assgn59012;
        z5901_assgn59014 <= z5901_assgn59013;
        z5901_assgn59015 <= z5901_assgn59014;
        z5901_assgn59016 <= z5901_assgn59015;
        z5901_assgn59017 <= z5901_assgn59016;
        z5901_assgn59018 <= z5901_assgn59017;
        z2125_assgn2125 <= z5901_assgn59018;
        z5913_assgn59130 <= z5913_assgn5913;
        z5913_assgn59131 <= z5913_assgn59130;
        z5913_assgn59132 <= z5913_assgn59131;
        z5913_assgn59133 <= z5913_assgn59132;
        z5913_assgn59134 <= z5913_assgn59133;
        z5913_assgn59135 <= z5913_assgn59134;
        z5913_assgn59136 <= z5913_assgn59135;
        z5913_assgn59137 <= z5913_assgn59136;
        z5913_assgn59138 <= z5913_assgn59137;
        z2135_assgn2135 <= z5913_assgn59138;
        z5917_assgn59170 <= z5917_assgn5917;
        z5917_assgn59171 <= z5917_assgn59170;
        z5917_assgn59172 <= z5917_assgn59171;
        z5917_assgn59173 <= z5917_assgn59172;
        z5917_assgn59174 <= z5917_assgn59173;
        z5917_assgn59175 <= z5917_assgn59174;
        z5917_assgn59176 <= z5917_assgn59175;
        z5917_assgn59177 <= z5917_assgn59176;
        z5917_assgn59178 <= z5917_assgn59177;
        z2137_assgn2137 <= z5917_assgn59178;
        z5925_assgn59250 <= z5925_assgn5925;
        z5925_assgn59251 <= z5925_assgn59250;
        z5925_assgn59252 <= z5925_assgn59251;
        z5925_assgn59253 <= z5925_assgn59252;
        z5925_assgn59254 <= z5925_assgn59253;
        z2143_assgn2143 <= z5925_assgn59254;
        z5929_assgn59290 <= z5929_assgn5929;
        z5929_assgn59291 <= z5929_assgn59290;
        z5929_assgn59292 <= z5929_assgn59291;
        z5929_assgn59293 <= z5929_assgn59292;
        z5929_assgn59294 <= z5929_assgn59293;
        z2145_assgn2145 <= z5929_assgn59294;
        z5933_assgn59330 <= z5933_assgn5933;
        z5933_assgn59331 <= z5933_assgn59330;
        z5933_assgn59332 <= z5933_assgn59331;
        z5933_assgn59333 <= z5933_assgn59332;
        z5933_assgn59334 <= z5933_assgn59333;
        z2147_assgn2147 <= z5933_assgn59334;
        z5937_assgn59370 <= z5937_assgn5937;
        z5937_assgn59371 <= z5937_assgn59370;
        z5937_assgn59372 <= z5937_assgn59371;
        z5937_assgn59373 <= z5937_assgn59372;
        z5937_assgn59374 <= z5937_assgn59373;
        z2149_assgn2149 <= z5937_assgn59374;
        z5941_assgn59410 <= z5941_assgn5941;
        z5941_assgn59411 <= z5941_assgn59410;
        z5941_assgn59412 <= z5941_assgn59411;
        z5941_assgn59413 <= z5941_assgn59412;
        z5941_assgn59414 <= z5941_assgn59413;
        z2151_assgn2151 <= z5941_assgn59414;
        z5945_assgn59450 <= z5945_assgn5945;
        z5945_assgn59451 <= z5945_assgn59450;
        z5945_assgn59452 <= z5945_assgn59451;
        z5945_assgn59453 <= z5945_assgn59452;
        z5945_assgn59454 <= z5945_assgn59453;
        z2153_assgn2153 <= z5945_assgn59454;
        z5949_assgn59490 <= z5949_assgn5949;
        z5949_assgn59491 <= z5949_assgn59490;
        z5949_assgn59492 <= z5949_assgn59491;
        z5949_assgn59493 <= z5949_assgn59492;
        z5949_assgn59494 <= z5949_assgn59493;
        z2155_assgn2155 <= z5949_assgn59494;
        z5953_assgn59530 <= z5953_assgn5953;
        z5953_assgn59531 <= z5953_assgn59530;
        z5953_assgn59532 <= z5953_assgn59531;
        z5953_assgn59533 <= z5953_assgn59532;
        z5953_assgn59534 <= z5953_assgn59533;
        z2157_assgn2157 <= z5953_assgn59534;
        z5957_assgn59570 <= z5957_assgn5957;
        z5957_assgn59571 <= z5957_assgn59570;
        z5957_assgn59572 <= z5957_assgn59571;
        z5957_assgn59573 <= z5957_assgn59572;
        z5957_assgn59574 <= z5957_assgn59573;
        z2159_assgn2159 <= z5957_assgn59574;
        z5961_assgn59610 <= z5961_assgn5961;
        z5961_assgn59611 <= z5961_assgn59610;
        z5961_assgn59612 <= z5961_assgn59611;
        z5961_assgn59613 <= z5961_assgn59612;
        z5961_assgn59614 <= z5961_assgn59613;
        z5961_assgn59615 <= z5961_assgn59614;
        z5961_assgn59616 <= z5961_assgn59615;
        z5961_assgn59617 <= z5961_assgn59616;
        z2161_assgn2161 <= z5961_assgn59617;
        z5965_assgn59650 <= z5965_assgn5965;
        z5965_assgn59651 <= z5965_assgn59650;
        z5965_assgn59652 <= z5965_assgn59651;
        z5965_assgn59653 <= z5965_assgn59652;
        z5965_assgn59654 <= z5965_assgn59653;
        z5965_assgn59655 <= z5965_assgn59654;
        z5965_assgn59656 <= z5965_assgn59655;
        z5965_assgn59657 <= z5965_assgn59656;
        z2163_assgn2163 <= z5965_assgn59657;
        z5969_assgn59690 <= z5969_assgn5969;
        z5969_assgn59691 <= z5969_assgn59690;
        z5969_assgn59692 <= z5969_assgn59691;
        z5969_assgn59693 <= z5969_assgn59692;
        z5969_assgn59694 <= z5969_assgn59693;
        z5969_assgn59695 <= z5969_assgn59694;
        z5969_assgn59696 <= z5969_assgn59695;
        z5969_assgn59697 <= z5969_assgn59696;
        z2165_assgn2165 <= z5969_assgn59697;
        z5973_assgn59730 <= z5973_assgn5973;
        z5973_assgn59731 <= z5973_assgn59730;
        z5973_assgn59732 <= z5973_assgn59731;
        z5973_assgn59733 <= z5973_assgn59732;
        z5973_assgn59734 <= z5973_assgn59733;
        z5973_assgn59735 <= z5973_assgn59734;
        z5973_assgn59736 <= z5973_assgn59735;
        z5973_assgn59737 <= z5973_assgn59736;
        z2167_assgn2167 <= z5973_assgn59737;
        z5977_assgn59770 <= z5977_assgn5977;
        z5977_assgn59771 <= z5977_assgn59770;
        z5977_assgn59772 <= z5977_assgn59771;
        z5977_assgn59773 <= z5977_assgn59772;
        z5977_assgn59774 <= z5977_assgn59773;
        z5977_assgn59775 <= z5977_assgn59774;
        z5977_assgn59776 <= z5977_assgn59775;
        z5977_assgn59777 <= z5977_assgn59776;
        z2169_assgn2169 <= z5977_assgn59777;
        z5981_assgn59810 <= z5981_assgn5981;
        z5981_assgn59811 <= z5981_assgn59810;
        z5981_assgn59812 <= z5981_assgn59811;
        z5981_assgn59813 <= z5981_assgn59812;
        z5981_assgn59814 <= z5981_assgn59813;
        z5981_assgn59815 <= z5981_assgn59814;
        z5981_assgn59816 <= z5981_assgn59815;
        z5981_assgn59817 <= z5981_assgn59816;
        z2171_assgn2171 <= z5981_assgn59817;
        z5985_assgn59850 <= z5985_assgn5985;
        z5985_assgn59851 <= z5985_assgn59850;
        z5985_assgn59852 <= z5985_assgn59851;
        z5985_assgn59853 <= z5985_assgn59852;
        z5985_assgn59854 <= z5985_assgn59853;
        z2173_assgn2173 <= z5985_assgn59854;
        z5987_assgn59870 <= z5987_assgn5987;
        z5987_assgn59871 <= z5987_assgn59870;
        z2174_assgn2174 <= z5987_assgn59871;
        z5991_assgn59910 <= z5991_assgn5991;
        z5991_assgn59911 <= z5991_assgn59910;
        z5991_assgn59912 <= z5991_assgn59911;
        z5991_assgn59913 <= z5991_assgn59912;
        z5991_assgn59914 <= z5991_assgn59913;
        z2175_assgn2175 <= z5991_assgn59914;
        z5993_assgn59930 <= z5993_assgn5993;
        z5993_assgn59931 <= z5993_assgn59930;
        z2176_assgn2176 <= z5993_assgn59931;
        z5997_assgn59970 <= z5997_assgn5997;
        z5997_assgn59971 <= z5997_assgn59970;
        z5997_assgn59972 <= z5997_assgn59971;
        z5997_assgn59973 <= z5997_assgn59972;
        z5997_assgn59974 <= z5997_assgn59973;
        z2177_assgn2177 <= z5997_assgn59974;
        z6001_assgn60010 <= z6001_assgn6001;
        z6001_assgn60011 <= z6001_assgn60010;
        z6001_assgn60012 <= z6001_assgn60011;
        z6001_assgn60013 <= z6001_assgn60012;
        z6001_assgn60014 <= z6001_assgn60013;
        z2179_assgn2179 <= z6001_assgn60014;
        z6005_assgn60050 <= z6005_assgn6005;
        z6005_assgn60051 <= z6005_assgn60050;
        z6005_assgn60052 <= z6005_assgn60051;
        z6005_assgn60053 <= z6005_assgn60052;
        z6005_assgn60054 <= z6005_assgn60053;
        z2181_assgn2181 <= z6005_assgn60054;
        z6007_assgn60070 <= z6007_assgn6007;
        z6007_assgn60071 <= z6007_assgn60070;
        z2182_assgn2182 <= z6007_assgn60071;
        z6011_assgn60110 <= z6011_assgn6011;
        z6011_assgn60111 <= z6011_assgn60110;
        z6011_assgn60112 <= z6011_assgn60111;
        z6011_assgn60113 <= z6011_assgn60112;
        z6011_assgn60114 <= z6011_assgn60113;
        z2183_assgn2183 <= z6011_assgn60114;
        z6013_assgn60130 <= z6013_assgn6013;
        z6013_assgn60131 <= z6013_assgn60130;
        z2184_assgn2184 <= z6013_assgn60131;
        z6025_assgn60250 <= z6025_assgn6025;
        z6025_assgn60251 <= z6025_assgn60250;
        z6025_assgn60252 <= z6025_assgn60251;
        z6025_assgn60253 <= z6025_assgn60252;
        z6025_assgn60254 <= z6025_assgn60253;
        z2193_assgn2193 <= z6025_assgn60254;
        z6029_assgn60290 <= z6029_assgn6029;
        z6029_assgn60291 <= z6029_assgn60290;
        z6029_assgn60292 <= z6029_assgn60291;
        z6029_assgn60293 <= z6029_assgn60292;
        z6029_assgn60294 <= z6029_assgn60293;
        z2195_assgn2195 <= z6029_assgn60294;
        z6033_assgn60330 <= z6033_assgn6033;
        z6033_assgn60331 <= z6033_assgn60330;
        z6033_assgn60332 <= z6033_assgn60331;
        z6033_assgn60333 <= z6033_assgn60332;
        z6033_assgn60334 <= z6033_assgn60333;
        z2197_assgn2197 <= z6033_assgn60334;
        z6037_assgn60370 <= z6037_assgn6037;
        z6037_assgn60371 <= z6037_assgn60370;
        z6037_assgn60372 <= z6037_assgn60371;
        z6037_assgn60373 <= z6037_assgn60372;
        z6037_assgn60374 <= z6037_assgn60373;
        z6037_assgn60375 <= z6037_assgn60374;
        z6037_assgn60376 <= z6037_assgn60375;
        z6037_assgn60377 <= z6037_assgn60376;
        z2199_assgn2199 <= z6037_assgn60377;
        z6041_assgn60410 <= z6041_assgn6041;
        z6041_assgn60411 <= z6041_assgn60410;
        z6041_assgn60412 <= z6041_assgn60411;
        z6041_assgn60413 <= z6041_assgn60412;
        z6041_assgn60414 <= z6041_assgn60413;
        z6041_assgn60415 <= z6041_assgn60414;
        z6041_assgn60416 <= z6041_assgn60415;
        z6041_assgn60417 <= z6041_assgn60416;
        z2201_assgn2201 <= z6041_assgn60417;
        z6045_assgn60450 <= z6045_assgn6045;
        z6045_assgn60451 <= z6045_assgn60450;
        z6045_assgn60452 <= z6045_assgn60451;
        z6045_assgn60453 <= z6045_assgn60452;
        z6045_assgn60454 <= z6045_assgn60453;
        z6045_assgn60455 <= z6045_assgn60454;
        z6045_assgn60456 <= z6045_assgn60455;
        z6045_assgn60457 <= z6045_assgn60456;
        z2203_assgn2203 <= z6045_assgn60457;
        z6049_assgn60490 <= z6049_assgn6049;
        z6049_assgn60491 <= z6049_assgn60490;
        z6049_assgn60492 <= z6049_assgn60491;
        z6049_assgn60493 <= z6049_assgn60492;
        z6049_assgn60494 <= z6049_assgn60493;
        z6049_assgn60495 <= z6049_assgn60494;
        z6049_assgn60496 <= z6049_assgn60495;
        z6049_assgn60497 <= z6049_assgn60496;
        z2205_assgn2205 <= z6049_assgn60497;
        z6053_assgn60530 <= z6053_assgn6053;
        z6053_assgn60531 <= z6053_assgn60530;
        z6053_assgn60532 <= z6053_assgn60531;
        z6053_assgn60533 <= z6053_assgn60532;
        z6053_assgn60534 <= z6053_assgn60533;
        z6053_assgn60535 <= z6053_assgn60534;
        z6053_assgn60536 <= z6053_assgn60535;
        z6053_assgn60537 <= z6053_assgn60536;
        z2207_assgn2207 <= z6053_assgn60537;
        z6057_assgn60570 <= z6057_assgn6057;
        z6057_assgn60571 <= z6057_assgn60570;
        z6057_assgn60572 <= z6057_assgn60571;
        z6057_assgn60573 <= z6057_assgn60572;
        z6057_assgn60574 <= z6057_assgn60573;
        z6057_assgn60575 <= z6057_assgn60574;
        z6057_assgn60576 <= z6057_assgn60575;
        z6057_assgn60577 <= z6057_assgn60576;
        z2209_assgn2209 <= z6057_assgn60577;
        z6061_assgn60610 <= z6061_assgn6061;
        z6061_assgn60611 <= z6061_assgn60610;
        z6061_assgn60612 <= z6061_assgn60611;
        z6061_assgn60613 <= z6061_assgn60612;
        z6061_assgn60614 <= z6061_assgn60613;
        z2211_assgn2211 <= z6061_assgn60614;
        z6065_assgn60650 <= z6065_assgn6065;
        z6065_assgn60651 <= z6065_assgn60650;
        z6065_assgn60652 <= z6065_assgn60651;
        z6065_assgn60653 <= z6065_assgn60652;
        z6065_assgn60654 <= z6065_assgn60653;
        z2213_assgn2213 <= z6065_assgn60654;
        z6069_assgn60690 <= z6069_assgn6069;
        z6069_assgn60691 <= z6069_assgn60690;
        z6069_assgn60692 <= z6069_assgn60691;
        z6069_assgn60693 <= z6069_assgn60692;
        z6069_assgn60694 <= z6069_assgn60693;
        z2215_assgn2215 <= z6069_assgn60694;
        z6073_assgn60730 <= z6073_assgn6073;
        z6073_assgn60731 <= z6073_assgn60730;
        z6073_assgn60732 <= z6073_assgn60731;
        z6073_assgn60733 <= z6073_assgn60732;
        z6073_assgn60734 <= z6073_assgn60733;
        z2217_assgn2217 <= z6073_assgn60734;
        z6077_assgn60770 <= z6077_assgn6077;
        z6077_assgn60771 <= z6077_assgn60770;
        z6077_assgn60772 <= z6077_assgn60771;
        z6077_assgn60773 <= z6077_assgn60772;
        z6077_assgn60774 <= z6077_assgn60773;
        z2219_assgn2219 <= z6077_assgn60774;
        z6081_assgn60810 <= z6081_assgn6081;
        z6081_assgn60811 <= z6081_assgn60810;
        z6081_assgn60812 <= z6081_assgn60811;
        z6081_assgn60813 <= z6081_assgn60812;
        z6081_assgn60814 <= z6081_assgn60813;
        z2221_assgn2221 <= z6081_assgn60814;
        c0_G4_mul0_G16_mul2_G256_inv0_reg <= c0_G4_mul0_G16_mul2_G256_inv0;
        d0_G4_mul0_G16_mul2_G256_inv0_reg <= d0_G4_mul0_G16_mul2_G256_inv0;
        c1_G4_mul0_G16_mul2_G256_inv0_reg <= c1_G4_mul0_G16_mul2_G256_inv0;
        d1_G4_mul0_G16_mul2_G256_inv0_reg <= d1_G4_mul0_G16_mul2_G256_inv0;
        z6093_assgn60930 <= z6093_assgn6093;
        z6093_assgn60931 <= z6093_assgn60930;
        z6093_assgn60932 <= z6093_assgn60931;
        z6093_assgn60933 <= z6093_assgn60932;
        z6093_assgn60934 <= z6093_assgn60933;
        z6093_assgn60935 <= z6093_assgn60934;
        z2231_assgn2231 <= z6093_assgn60935;
        z6101_assgn61010 <= z6101_assgn6101;
        z2237_assgn2237 <= z6101_assgn61010;
        z6105_assgn61050 <= z6105_assgn6105;
        z2239_assgn2239 <= z6105_assgn61050;
        cxord_0_G4_mul0_G16_mul2_G256_inv0_reg <= cxord_0_G4_mul0_G16_mul2_G256_inv0;
        r0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
        cxord_1_G4_mul0_G16_mul2_G256_inv0_reg <= cxord_1_G4_mul0_G16_mul2_G256_inv0;
        z6113_assgn61130 <= z6113_assgn6113;
        z2245_assgn2245 <= z6113_assgn61130;
        v1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= v1_hpc20_G4_mul0_G16_mul2_G256_inv0;
        u0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= u0_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p0_hpc20_G4_mul0_G16_mul2_G256_inv0;
        z6123_assgn61230 <= z6123_assgn6123;
        z2253_assgn2253 <= z6123_assgn61230;
        v0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= v0_hpc20_G4_mul0_G16_mul2_G256_inv0;
        u1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= u1_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p3_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p3_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p2_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p2_hpc20_G4_mul0_G16_mul2_G256_inv0;
        z6133_assgn61330 <= z6133_assgn6133;
        z6133_assgn61331 <= z6133_assgn61330;
        z6133_assgn61332 <= z6133_assgn61331;
        z6133_assgn61333 <= z6133_assgn61332;
        z6133_assgn61334 <= z6133_assgn61333;
        z6133_assgn61335 <= z6133_assgn61334;
        z2261_assgn2261 <= z6133_assgn61335;
        z6141_assgn61410 <= z6141_assgn6141;
        z2267_assgn2267 <= z6141_assgn61410;
        z6145_assgn61450 <= z6145_assgn6145;
        z2269_assgn2269 <= z6145_assgn61450;
        z6149_assgn61490 <= z6149_assgn6149;
        z2272_assgn2272 <= z6149_assgn61490;
        r0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
        z6153_assgn61530 <= z6153_assgn6153;
        z2274_assgn2274 <= z6153_assgn61530;
        z6157_assgn61570 <= z6157_assgn6157;
        z6157_assgn61571 <= z6157_assgn61570;
        z2275_assgn2275 <= z6157_assgn61571;
        v1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= v1_hpc21_G4_mul0_G16_mul2_G256_inv0;
        u0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= u0_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p0_hpc21_G4_mul0_G16_mul2_G256_inv0;
        z6167_assgn61670 <= z6167_assgn6167;
        z6167_assgn61671 <= z6167_assgn61670;
        z2283_assgn2283 <= z6167_assgn61671;
        v0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= v0_hpc21_G4_mul0_G16_mul2_G256_inv0;
        u1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= u1_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p3_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p3_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p2_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p2_hpc21_G4_mul0_G16_mul2_G256_inv0;
        z6181_assgn61810 <= z6181_assgn6181;
        z6181_assgn61811 <= z6181_assgn61810;
        z6181_assgn61812 <= z6181_assgn61811;
        z6181_assgn61813 <= z6181_assgn61812;
        z6181_assgn61814 <= z6181_assgn61813;
        z6181_assgn61815 <= z6181_assgn61814;
        z2295_assgn2295 <= z6181_assgn61815;
        z6189_assgn61890 <= z6189_assgn6189;
        z2301_assgn2301 <= z6189_assgn61890;
        z6193_assgn61930 <= z6193_assgn6193;
        z2303_assgn2303 <= z6193_assgn61930;
        z6197_assgn61970 <= z6197_assgn6197;
        z2306_assgn2306 <= z6197_assgn61970;
        r0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
        z6201_assgn62010 <= z6201_assgn6201;
        z2308_assgn2308 <= z6201_assgn62010;
        z6205_assgn62050 <= z6205_assgn6205;
        z6205_assgn62051 <= z6205_assgn62050;
        z2309_assgn2309 <= z6205_assgn62051;
        v1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= v1_hpc22_G4_mul0_G16_mul2_G256_inv0;
        u0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= u0_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p0_hpc22_G4_mul0_G16_mul2_G256_inv0;
        z6215_assgn62150 <= z6215_assgn6215;
        z6215_assgn62151 <= z6215_assgn62150;
        z2317_assgn2317 <= z6215_assgn62151;
        v0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= v0_hpc22_G4_mul0_G16_mul2_G256_inv0;
        u1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= u1_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p3_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p3_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p2_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p2_hpc22_G4_mul0_G16_mul2_G256_inv0;
        z6229_assgn62290 <= z6229_assgn6229;
        z6229_assgn62291 <= z6229_assgn62290;
        z6229_assgn62292 <= z6229_assgn62291;
        z6229_assgn62293 <= z6229_assgn62292;
        z6229_assgn62294 <= z6229_assgn62293;
        z6229_assgn62295 <= z6229_assgn62294;
        z6229_assgn62296 <= z6229_assgn62295;
        z6229_assgn62297 <= z6229_assgn62296;
        z6229_assgn62298 <= z6229_assgn62297;
        z2329_assgn2329 <= z6229_assgn62298;
        z6233_assgn62330 <= z6233_assgn6233;
        z6233_assgn62331 <= z6233_assgn62330;
        z6233_assgn62332 <= z6233_assgn62331;
        z6233_assgn62333 <= z6233_assgn62332;
        z6233_assgn62334 <= z6233_assgn62333;
        z6233_assgn62335 <= z6233_assgn62334;
        z6233_assgn62336 <= z6233_assgn62335;
        z6233_assgn62337 <= z6233_assgn62336;
        z6233_assgn62338 <= z6233_assgn62337;
        z2331_assgn2331 <= z6233_assgn62338;
        z6241_assgn62410 <= z6241_assgn6241;
        z6241_assgn62411 <= z6241_assgn62410;
        z6241_assgn62412 <= z6241_assgn62411;
        z6241_assgn62413 <= z6241_assgn62412;
        z6241_assgn62414 <= z6241_assgn62413;
        z6241_assgn62415 <= z6241_assgn62414;
        z6241_assgn62416 <= z6241_assgn62415;
        z6241_assgn62417 <= z6241_assgn62416;
        z6241_assgn62418 <= z6241_assgn62417;
        z2337_assgn2337 <= z6241_assgn62418;
        z6245_assgn62450 <= z6245_assgn6245;
        z6245_assgn62451 <= z6245_assgn62450;
        z6245_assgn62452 <= z6245_assgn62451;
        z6245_assgn62453 <= z6245_assgn62452;
        z6245_assgn62454 <= z6245_assgn62453;
        z6245_assgn62455 <= z6245_assgn62454;
        z6245_assgn62456 <= z6245_assgn62455;
        z6245_assgn62457 <= z6245_assgn62456;
        z6245_assgn62458 <= z6245_assgn62457;
        z2339_assgn2339 <= z6245_assgn62458;
        z6249_assgn62490 <= z6249_assgn6249;
        z6249_assgn62491 <= z6249_assgn62490;
        z6249_assgn62492 <= z6249_assgn62491;
        z6249_assgn62493 <= z6249_assgn62492;
        z6249_assgn62494 <= z6249_assgn62493;
        z6249_assgn62495 <= z6249_assgn62494;
        z6249_assgn62496 <= z6249_assgn62495;
        z6249_assgn62497 <= z6249_assgn62496;
        z6249_assgn62498 <= z6249_assgn62497;
        z2341_assgn2341 <= z6249_assgn62498;
        z6253_assgn62530 <= z6253_assgn6253;
        z6253_assgn62531 <= z6253_assgn62530;
        z6253_assgn62532 <= z6253_assgn62531;
        z6253_assgn62533 <= z6253_assgn62532;
        z6253_assgn62534 <= z6253_assgn62533;
        z6253_assgn62535 <= z6253_assgn62534;
        z6253_assgn62536 <= z6253_assgn62535;
        z6253_assgn62537 <= z6253_assgn62536;
        z6253_assgn62538 <= z6253_assgn62537;
        z2343_assgn2343 <= z6253_assgn62538;
        z6257_assgn62570 <= z6257_assgn6257;
        z6257_assgn62571 <= z6257_assgn62570;
        z6257_assgn62572 <= z6257_assgn62571;
        z6257_assgn62573 <= z6257_assgn62572;
        z6257_assgn62574 <= z6257_assgn62573;
        z6257_assgn62575 <= z6257_assgn62574;
        z6257_assgn62576 <= z6257_assgn62575;
        z6257_assgn62577 <= z6257_assgn62576;
        z6257_assgn62578 <= z6257_assgn62577;
        z2345_assgn2345 <= z6257_assgn62578;
        z6261_assgn62610 <= z6261_assgn6261;
        z6261_assgn62611 <= z6261_assgn62610;
        z6261_assgn62612 <= z6261_assgn62611;
        z6261_assgn62613 <= z6261_assgn62612;
        z6261_assgn62614 <= z6261_assgn62613;
        z6261_assgn62615 <= z6261_assgn62614;
        z6261_assgn62616 <= z6261_assgn62615;
        z6261_assgn62617 <= z6261_assgn62616;
        z6261_assgn62618 <= z6261_assgn62617;
        z2347_assgn2347 <= z6261_assgn62618;
        z6273_assgn62730 <= z6273_assgn6273;
        z6273_assgn62731 <= z6273_assgn62730;
        z6273_assgn62732 <= z6273_assgn62731;
        z6273_assgn62733 <= z6273_assgn62732;
        z6273_assgn62734 <= z6273_assgn62733;
        z6273_assgn62735 <= z6273_assgn62734;
        z6273_assgn62736 <= z6273_assgn62735;
        z6273_assgn62737 <= z6273_assgn62736;
        z6273_assgn62738 <= z6273_assgn62737;
        z2357_assgn2357 <= z6273_assgn62738;
        z6277_assgn62770 <= z6277_assgn6277;
        z6277_assgn62771 <= z6277_assgn62770;
        z6277_assgn62772 <= z6277_assgn62771;
        z6277_assgn62773 <= z6277_assgn62772;
        z6277_assgn62774 <= z6277_assgn62773;
        z6277_assgn62775 <= z6277_assgn62774;
        z6277_assgn62776 <= z6277_assgn62775;
        z6277_assgn62777 <= z6277_assgn62776;
        z6277_assgn62778 <= z6277_assgn62777;
        z2359_assgn2359 <= z6277_assgn62778;
        z6285_assgn62850 <= z6285_assgn6285;
        z6285_assgn62851 <= z6285_assgn62850;
        z6285_assgn62852 <= z6285_assgn62851;
        z6285_assgn62853 <= z6285_assgn62852;
        z6285_assgn62854 <= z6285_assgn62853;
        z2365_assgn2365 <= z6285_assgn62854;
        z6289_assgn62890 <= z6289_assgn6289;
        z6289_assgn62891 <= z6289_assgn62890;
        z6289_assgn62892 <= z6289_assgn62891;
        z6289_assgn62893 <= z6289_assgn62892;
        z6289_assgn62894 <= z6289_assgn62893;
        z2367_assgn2367 <= z6289_assgn62894;
        z6293_assgn62930 <= z6293_assgn6293;
        z6293_assgn62931 <= z6293_assgn62930;
        z6293_assgn62932 <= z6293_assgn62931;
        z6293_assgn62933 <= z6293_assgn62932;
        z6293_assgn62934 <= z6293_assgn62933;
        z2369_assgn2369 <= z6293_assgn62934;
        z6297_assgn62970 <= z6297_assgn6297;
        z6297_assgn62971 <= z6297_assgn62970;
        z6297_assgn62972 <= z6297_assgn62971;
        z6297_assgn62973 <= z6297_assgn62972;
        z6297_assgn62974 <= z6297_assgn62973;
        z6297_assgn62975 <= z6297_assgn62974;
        z6297_assgn62976 <= z6297_assgn62975;
        z6297_assgn62977 <= z6297_assgn62976;
        z2371_assgn2371 <= z6297_assgn62977;
        z6301_assgn63010 <= z6301_assgn6301;
        z6301_assgn63011 <= z6301_assgn63010;
        z6301_assgn63012 <= z6301_assgn63011;
        z6301_assgn63013 <= z6301_assgn63012;
        z6301_assgn63014 <= z6301_assgn63013;
        z6301_assgn63015 <= z6301_assgn63014;
        z6301_assgn63016 <= z6301_assgn63015;
        z6301_assgn63017 <= z6301_assgn63016;
        z2373_assgn2373 <= z6301_assgn63017;
        z6305_assgn63050 <= z6305_assgn6305;
        z6305_assgn63051 <= z6305_assgn63050;
        z6305_assgn63052 <= z6305_assgn63051;
        z6305_assgn63053 <= z6305_assgn63052;
        z6305_assgn63054 <= z6305_assgn63053;
        z6305_assgn63055 <= z6305_assgn63054;
        z6305_assgn63056 <= z6305_assgn63055;
        z6305_assgn63057 <= z6305_assgn63056;
        z2375_assgn2375 <= z6305_assgn63057;
        z6309_assgn63090 <= z6309_assgn6309;
        z6309_assgn63091 <= z6309_assgn63090;
        z6309_assgn63092 <= z6309_assgn63091;
        z6309_assgn63093 <= z6309_assgn63092;
        z6309_assgn63094 <= z6309_assgn63093;
        z6309_assgn63095 <= z6309_assgn63094;
        z6309_assgn63096 <= z6309_assgn63095;
        z6309_assgn63097 <= z6309_assgn63096;
        z2377_assgn2377 <= z6309_assgn63097;
        z6313_assgn63130 <= z6313_assgn6313;
        z6313_assgn63131 <= z6313_assgn63130;
        z6313_assgn63132 <= z6313_assgn63131;
        z6313_assgn63133 <= z6313_assgn63132;
        z6313_assgn63134 <= z6313_assgn63133;
        z6313_assgn63135 <= z6313_assgn63134;
        z6313_assgn63136 <= z6313_assgn63135;
        z6313_assgn63137 <= z6313_assgn63136;
        z2379_assgn2379 <= z6313_assgn63137;
        z6317_assgn63170 <= z6317_assgn6317;
        z6317_assgn63171 <= z6317_assgn63170;
        z6317_assgn63172 <= z6317_assgn63171;
        z6317_assgn63173 <= z6317_assgn63172;
        z6317_assgn63174 <= z6317_assgn63173;
        z6317_assgn63175 <= z6317_assgn63174;
        z6317_assgn63176 <= z6317_assgn63175;
        z6317_assgn63177 <= z6317_assgn63176;
        z2381_assgn2381 <= z6317_assgn63177;
        z6321_assgn63210 <= z6321_assgn6321;
        z6321_assgn63211 <= z6321_assgn63210;
        z6321_assgn63212 <= z6321_assgn63211;
        z6321_assgn63213 <= z6321_assgn63212;
        z6321_assgn63214 <= z6321_assgn63213;
        z2383_assgn2383 <= z6321_assgn63214;
        z6325_assgn63250 <= z6325_assgn6325;
        z6325_assgn63251 <= z6325_assgn63250;
        z6325_assgn63252 <= z6325_assgn63251;
        z6325_assgn63253 <= z6325_assgn63252;
        z6325_assgn63254 <= z6325_assgn63253;
        z2385_assgn2385 <= z6325_assgn63254;
        z6329_assgn63290 <= z6329_assgn6329;
        z6329_assgn63291 <= z6329_assgn63290;
        z6329_assgn63292 <= z6329_assgn63291;
        z6329_assgn63293 <= z6329_assgn63292;
        z6329_assgn63294 <= z6329_assgn63293;
        z2387_assgn2387 <= z6329_assgn63294;
        z6333_assgn63330 <= z6333_assgn6333;
        z6333_assgn63331 <= z6333_assgn63330;
        z6333_assgn63332 <= z6333_assgn63331;
        z6333_assgn63333 <= z6333_assgn63332;
        z6333_assgn63334 <= z6333_assgn63333;
        z2389_assgn2389 <= z6333_assgn63334;
        z6337_assgn63370 <= z6337_assgn6337;
        z6337_assgn63371 <= z6337_assgn63370;
        z6337_assgn63372 <= z6337_assgn63371;
        z6337_assgn63373 <= z6337_assgn63372;
        z6337_assgn63374 <= z6337_assgn63373;
        z2391_assgn2391 <= z6337_assgn63374;
        z6341_assgn63410 <= z6341_assgn6341;
        z6341_assgn63411 <= z6341_assgn63410;
        z6341_assgn63412 <= z6341_assgn63411;
        z6341_assgn63413 <= z6341_assgn63412;
        z6341_assgn63414 <= z6341_assgn63413;
        z2393_assgn2393 <= z6341_assgn63414;
        c0_G4_mul1_G16_mul2_G256_inv0_reg <= c0_G4_mul1_G16_mul2_G256_inv0;
        d0_G4_mul1_G16_mul2_G256_inv0_reg <= d0_G4_mul1_G16_mul2_G256_inv0;
        c1_G4_mul1_G16_mul2_G256_inv0_reg <= c1_G4_mul1_G16_mul2_G256_inv0;
        d1_G4_mul1_G16_mul2_G256_inv0_reg <= d1_G4_mul1_G16_mul2_G256_inv0;
        z6353_assgn63530 <= z6353_assgn6353;
        z6353_assgn63531 <= z6353_assgn63530;
        z6353_assgn63532 <= z6353_assgn63531;
        z6353_assgn63533 <= z6353_assgn63532;
        z6353_assgn63534 <= z6353_assgn63533;
        z6353_assgn63535 <= z6353_assgn63534;
        z2403_assgn2403 <= z6353_assgn63535;
        z6361_assgn63610 <= z6361_assgn6361;
        z2409_assgn2409 <= z6361_assgn63610;
        z6365_assgn63650 <= z6365_assgn6365;
        z2411_assgn2411 <= z6365_assgn63650;
        cxord_0_G4_mul1_G16_mul2_G256_inv0_reg <= cxord_0_G4_mul1_G16_mul2_G256_inv0;
        r0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
        cxord_1_G4_mul1_G16_mul2_G256_inv0_reg <= cxord_1_G4_mul1_G16_mul2_G256_inv0;
        z6373_assgn63730 <= z6373_assgn6373;
        z2417_assgn2417 <= z6373_assgn63730;
        v1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= v1_hpc20_G4_mul1_G16_mul2_G256_inv0;
        u0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= u0_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p0_hpc20_G4_mul1_G16_mul2_G256_inv0;
        z6383_assgn63830 <= z6383_assgn6383;
        z2425_assgn2425 <= z6383_assgn63830;
        v0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= v0_hpc20_G4_mul1_G16_mul2_G256_inv0;
        u1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= u1_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p3_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p3_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p2_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p2_hpc20_G4_mul1_G16_mul2_G256_inv0;
        z6393_assgn63930 <= z6393_assgn6393;
        z6393_assgn63931 <= z6393_assgn63930;
        z6393_assgn63932 <= z6393_assgn63931;
        z6393_assgn63933 <= z6393_assgn63932;
        z6393_assgn63934 <= z6393_assgn63933;
        z6393_assgn63935 <= z6393_assgn63934;
        z2433_assgn2433 <= z6393_assgn63935;
        z6401_assgn64010 <= z6401_assgn6401;
        z2439_assgn2439 <= z6401_assgn64010;
        z6405_assgn64050 <= z6405_assgn6405;
        z2441_assgn2441 <= z6405_assgn64050;
        z6409_assgn64090 <= z6409_assgn6409;
        z2444_assgn2444 <= z6409_assgn64090;
        r0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
        z6413_assgn64130 <= z6413_assgn6413;
        z2446_assgn2446 <= z6413_assgn64130;
        z6417_assgn64170 <= z6417_assgn6417;
        z6417_assgn64171 <= z6417_assgn64170;
        z2447_assgn2447 <= z6417_assgn64171;
        v1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= v1_hpc21_G4_mul1_G16_mul2_G256_inv0;
        u0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= u0_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p0_hpc21_G4_mul1_G16_mul2_G256_inv0;
        z6427_assgn64270 <= z6427_assgn6427;
        z6427_assgn64271 <= z6427_assgn64270;
        z2455_assgn2455 <= z6427_assgn64271;
        v0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= v0_hpc21_G4_mul1_G16_mul2_G256_inv0;
        u1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= u1_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p3_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p3_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p2_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p2_hpc21_G4_mul1_G16_mul2_G256_inv0;
        z6441_assgn64410 <= z6441_assgn6441;
        z6441_assgn64411 <= z6441_assgn64410;
        z6441_assgn64412 <= z6441_assgn64411;
        z6441_assgn64413 <= z6441_assgn64412;
        z6441_assgn64414 <= z6441_assgn64413;
        z6441_assgn64415 <= z6441_assgn64414;
        z2467_assgn2467 <= z6441_assgn64415;
        z6449_assgn64490 <= z6449_assgn6449;
        z2473_assgn2473 <= z6449_assgn64490;
        z6453_assgn64530 <= z6453_assgn6453;
        z2475_assgn2475 <= z6453_assgn64530;
        z6457_assgn64570 <= z6457_assgn6457;
        z2478_assgn2478 <= z6457_assgn64570;
        r0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
        z6461_assgn64610 <= z6461_assgn6461;
        z2480_assgn2480 <= z6461_assgn64610;
        z6465_assgn64650 <= z6465_assgn6465;
        z6465_assgn64651 <= z6465_assgn64650;
        z2481_assgn2481 <= z6465_assgn64651;
        v1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= v1_hpc22_G4_mul1_G16_mul2_G256_inv0;
        u0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= u0_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p0_hpc22_G4_mul1_G16_mul2_G256_inv0;
        z6475_assgn64750 <= z6475_assgn6475;
        z6475_assgn64751 <= z6475_assgn64750;
        z2489_assgn2489 <= z6475_assgn64751;
        v0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= v0_hpc22_G4_mul1_G16_mul2_G256_inv0;
        u1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= u1_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p3_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p3_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p2_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p2_hpc22_G4_mul1_G16_mul2_G256_inv0;
        z6489_assgn64890 <= z6489_assgn6489;
        z6489_assgn64891 <= z6489_assgn64890;
        z6489_assgn64892 <= z6489_assgn64891;
        z6489_assgn64893 <= z6489_assgn64892;
        z6489_assgn64894 <= z6489_assgn64893;
        z6489_assgn64895 <= z6489_assgn64894;
        z6489_assgn64896 <= z6489_assgn64895;
        z6489_assgn64897 <= z6489_assgn64896;
        z6489_assgn64898 <= z6489_assgn64897;
        z2501_assgn2501 <= z6489_assgn64898;
        z6493_assgn64930 <= z6493_assgn6493;
        z6493_assgn64931 <= z6493_assgn64930;
        z6493_assgn64932 <= z6493_assgn64931;
        z6493_assgn64933 <= z6493_assgn64932;
        z6493_assgn64934 <= z6493_assgn64933;
        z6493_assgn64935 <= z6493_assgn64934;
        z6493_assgn64936 <= z6493_assgn64935;
        z6493_assgn64937 <= z6493_assgn64936;
        z6493_assgn64938 <= z6493_assgn64937;
        z2503_assgn2503 <= z6493_assgn64938;
        z6505_assgn65050 <= z6505_assgn6505;
        z6505_assgn65051 <= z6505_assgn65050;
        z6505_assgn65052 <= z6505_assgn65051;
        z6505_assgn65053 <= z6505_assgn65052;
        z6505_assgn65054 <= z6505_assgn65053;
        z2513_assgn2513 <= z6505_assgn65054;
        z6509_assgn65090 <= z6509_assgn6509;
        z6509_assgn65091 <= z6509_assgn65090;
        z6509_assgn65092 <= z6509_assgn65091;
        z6509_assgn65093 <= z6509_assgn65092;
        z6509_assgn65094 <= z6509_assgn65093;
        z2515_assgn2515 <= z6509_assgn65094;
        z6513_assgn65130 <= z6513_assgn6513;
        z6513_assgn65131 <= z6513_assgn65130;
        z6513_assgn65132 <= z6513_assgn65131;
        z6513_assgn65133 <= z6513_assgn65132;
        z6513_assgn65134 <= z6513_assgn65133;
        z2517_assgn2517 <= z6513_assgn65134;
        z6517_assgn65170 <= z6517_assgn6517;
        z6517_assgn65171 <= z6517_assgn65170;
        z6517_assgn65172 <= z6517_assgn65171;
        z6517_assgn65173 <= z6517_assgn65172;
        z6517_assgn65174 <= z6517_assgn65173;
        z6517_assgn65175 <= z6517_assgn65174;
        z6517_assgn65176 <= z6517_assgn65175;
        z6517_assgn65177 <= z6517_assgn65176;
        z2519_assgn2519 <= z6517_assgn65177;
        z6521_assgn65210 <= z6521_assgn6521;
        z6521_assgn65211 <= z6521_assgn65210;
        z6521_assgn65212 <= z6521_assgn65211;
        z6521_assgn65213 <= z6521_assgn65212;
        z6521_assgn65214 <= z6521_assgn65213;
        z6521_assgn65215 <= z6521_assgn65214;
        z6521_assgn65216 <= z6521_assgn65215;
        z6521_assgn65217 <= z6521_assgn65216;
        z2521_assgn2521 <= z6521_assgn65217;
        z6525_assgn65250 <= z6525_assgn6525;
        z6525_assgn65251 <= z6525_assgn65250;
        z6525_assgn65252 <= z6525_assgn65251;
        z6525_assgn65253 <= z6525_assgn65252;
        z6525_assgn65254 <= z6525_assgn65253;
        z6525_assgn65255 <= z6525_assgn65254;
        z6525_assgn65256 <= z6525_assgn65255;
        z6525_assgn65257 <= z6525_assgn65256;
        z2523_assgn2523 <= z6525_assgn65257;
        z6529_assgn65290 <= z6529_assgn6529;
        z6529_assgn65291 <= z6529_assgn65290;
        z6529_assgn65292 <= z6529_assgn65291;
        z6529_assgn65293 <= z6529_assgn65292;
        z6529_assgn65294 <= z6529_assgn65293;
        z6529_assgn65295 <= z6529_assgn65294;
        z6529_assgn65296 <= z6529_assgn65295;
        z6529_assgn65297 <= z6529_assgn65296;
        z2525_assgn2525 <= z6529_assgn65297;
        z6533_assgn65330 <= z6533_assgn6533;
        z6533_assgn65331 <= z6533_assgn65330;
        z6533_assgn65332 <= z6533_assgn65331;
        z6533_assgn65333 <= z6533_assgn65332;
        z6533_assgn65334 <= z6533_assgn65333;
        z6533_assgn65335 <= z6533_assgn65334;
        z6533_assgn65336 <= z6533_assgn65335;
        z6533_assgn65337 <= z6533_assgn65336;
        z2527_assgn2527 <= z6533_assgn65337;
        z6537_assgn65370 <= z6537_assgn6537;
        z6537_assgn65371 <= z6537_assgn65370;
        z6537_assgn65372 <= z6537_assgn65371;
        z6537_assgn65373 <= z6537_assgn65372;
        z6537_assgn65374 <= z6537_assgn65373;
        z6537_assgn65375 <= z6537_assgn65374;
        z6537_assgn65376 <= z6537_assgn65375;
        z6537_assgn65377 <= z6537_assgn65376;
        z2529_assgn2529 <= z6537_assgn65377;
        z6541_assgn65410 <= z6541_assgn6541;
        z6541_assgn65411 <= z6541_assgn65410;
        z6541_assgn65412 <= z6541_assgn65411;
        z6541_assgn65413 <= z6541_assgn65412;
        z6541_assgn65414 <= z6541_assgn65413;
        z2531_assgn2531 <= z6541_assgn65414;
        z6545_assgn65450 <= z6545_assgn6545;
        z6545_assgn65451 <= z6545_assgn65450;
        z6545_assgn65452 <= z6545_assgn65451;
        z6545_assgn65453 <= z6545_assgn65452;
        z6545_assgn65454 <= z6545_assgn65453;
        z2533_assgn2533 <= z6545_assgn65454;
        z6549_assgn65490 <= z6549_assgn6549;
        z6549_assgn65491 <= z6549_assgn65490;
        z6549_assgn65492 <= z6549_assgn65491;
        z6549_assgn65493 <= z6549_assgn65492;
        z6549_assgn65494 <= z6549_assgn65493;
        z2535_assgn2535 <= z6549_assgn65494;
        z6553_assgn65530 <= z6553_assgn6553;
        z6553_assgn65531 <= z6553_assgn65530;
        z6553_assgn65532 <= z6553_assgn65531;
        z6553_assgn65533 <= z6553_assgn65532;
        z6553_assgn65534 <= z6553_assgn65533;
        z2537_assgn2537 <= z6553_assgn65534;
        z6557_assgn65570 <= z6557_assgn6557;
        z6557_assgn65571 <= z6557_assgn65570;
        z6557_assgn65572 <= z6557_assgn65571;
        z6557_assgn65573 <= z6557_assgn65572;
        z6557_assgn65574 <= z6557_assgn65573;
        z2539_assgn2539 <= z6557_assgn65574;
        z6561_assgn65610 <= z6561_assgn6561;
        z6561_assgn65611 <= z6561_assgn65610;
        z6561_assgn65612 <= z6561_assgn65611;
        z6561_assgn65613 <= z6561_assgn65612;
        z6561_assgn65614 <= z6561_assgn65613;
        z2541_assgn2541 <= z6561_assgn65614;
        c0_G4_mul2_G16_mul2_G256_inv0_reg <= c0_G4_mul2_G16_mul2_G256_inv0;
        d0_G4_mul2_G16_mul2_G256_inv0_reg <= d0_G4_mul2_G16_mul2_G256_inv0;
        c1_G4_mul2_G16_mul2_G256_inv0_reg <= c1_G4_mul2_G16_mul2_G256_inv0;
        d1_G4_mul2_G16_mul2_G256_inv0_reg <= d1_G4_mul2_G16_mul2_G256_inv0;
        z6573_assgn65730 <= z6573_assgn6573;
        z6573_assgn65731 <= z6573_assgn65730;
        z6573_assgn65732 <= z6573_assgn65731;
        z6573_assgn65733 <= z6573_assgn65732;
        z6573_assgn65734 <= z6573_assgn65733;
        z6573_assgn65735 <= z6573_assgn65734;
        z2551_assgn2551 <= z6573_assgn65735;
        z6581_assgn65810 <= z6581_assgn6581;
        z2557_assgn2557 <= z6581_assgn65810;
        z6585_assgn65850 <= z6585_assgn6585;
        z2559_assgn2559 <= z6585_assgn65850;
        cxord_0_G4_mul2_G16_mul2_G256_inv0_reg <= cxord_0_G4_mul2_G16_mul2_G256_inv0;
        r0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
        cxord_1_G4_mul2_G16_mul2_G256_inv0_reg <= cxord_1_G4_mul2_G16_mul2_G256_inv0;
        z6593_assgn65930 <= z6593_assgn6593;
        z2565_assgn2565 <= z6593_assgn65930;
        v1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= v1_hpc20_G4_mul2_G16_mul2_G256_inv0;
        u0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= u0_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p0_hpc20_G4_mul2_G16_mul2_G256_inv0;
        z6603_assgn66030 <= z6603_assgn6603;
        z2573_assgn2573 <= z6603_assgn66030;
        v0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= v0_hpc20_G4_mul2_G16_mul2_G256_inv0;
        u1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= u1_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p3_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p3_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p2_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p2_hpc20_G4_mul2_G16_mul2_G256_inv0;
        z6613_assgn66130 <= z6613_assgn6613;
        z6613_assgn66131 <= z6613_assgn66130;
        z6613_assgn66132 <= z6613_assgn66131;
        z6613_assgn66133 <= z6613_assgn66132;
        z6613_assgn66134 <= z6613_assgn66133;
        z6613_assgn66135 <= z6613_assgn66134;
        z2581_assgn2581 <= z6613_assgn66135;
        z6621_assgn66210 <= z6621_assgn6621;
        z2587_assgn2587 <= z6621_assgn66210;
        z6625_assgn66250 <= z6625_assgn6625;
        z2589_assgn2589 <= z6625_assgn66250;
        z6629_assgn66290 <= z6629_assgn6629;
        z2592_assgn2592 <= z6629_assgn66290;
        r0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
        z6633_assgn66330 <= z6633_assgn6633;
        z2594_assgn2594 <= z6633_assgn66330;
        z6637_assgn66370 <= z6637_assgn6637;
        z6637_assgn66371 <= z6637_assgn66370;
        z2595_assgn2595 <= z6637_assgn66371;
        v1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= v1_hpc21_G4_mul2_G16_mul2_G256_inv0;
        u0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= u0_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p0_hpc21_G4_mul2_G16_mul2_G256_inv0;
        z6647_assgn66470 <= z6647_assgn6647;
        z6647_assgn66471 <= z6647_assgn66470;
        z2603_assgn2603 <= z6647_assgn66471;
        v0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= v0_hpc21_G4_mul2_G16_mul2_G256_inv0;
        u1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= u1_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p3_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p3_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p2_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p2_hpc21_G4_mul2_G16_mul2_G256_inv0;
        z6661_assgn66610 <= z6661_assgn6661;
        z6661_assgn66611 <= z6661_assgn66610;
        z6661_assgn66612 <= z6661_assgn66611;
        z6661_assgn66613 <= z6661_assgn66612;
        z6661_assgn66614 <= z6661_assgn66613;
        z6661_assgn66615 <= z6661_assgn66614;
        z2615_assgn2615 <= z6661_assgn66615;
        z6669_assgn66690 <= z6669_assgn6669;
        z2621_assgn2621 <= z6669_assgn66690;
        z6673_assgn66730 <= z6673_assgn6673;
        z2623_assgn2623 <= z6673_assgn66730;
        z6677_assgn66770 <= z6677_assgn6677;
        z2626_assgn2626 <= z6677_assgn66770;
        r0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
        z6681_assgn66810 <= z6681_assgn6681;
        z2628_assgn2628 <= z6681_assgn66810;
        z6685_assgn66850 <= z6685_assgn6685;
        z6685_assgn66851 <= z6685_assgn66850;
        z2629_assgn2629 <= z6685_assgn66851;
        v1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= v1_hpc22_G4_mul2_G16_mul2_G256_inv0;
        u0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= u0_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p0_hpc22_G4_mul2_G16_mul2_G256_inv0;
        z6695_assgn66950 <= z6695_assgn6695;
        z6695_assgn66951 <= z6695_assgn66950;
        z2637_assgn2637 <= z6695_assgn66951;
        v0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= v0_hpc22_G4_mul2_G16_mul2_G256_inv0;
        u1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= u1_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p3_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p3_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p2_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p2_hpc22_G4_mul2_G16_mul2_G256_inv0;
        z6709_assgn67090 <= z6709_assgn6709;
        z6709_assgn67091 <= z6709_assgn67090;
        z6709_assgn67092 <= z6709_assgn67091;
        z6709_assgn67093 <= z6709_assgn67092;
        z6709_assgn67094 <= z6709_assgn67093;
        z6709_assgn67095 <= z6709_assgn67094;
        z6709_assgn67096 <= z6709_assgn67095;
        z6709_assgn67097 <= z6709_assgn67096;
        z6709_assgn67098 <= z6709_assgn67097;
        z2649_assgn2649 <= z6709_assgn67098;
        z6713_assgn67130 <= z6713_assgn6713;
        z6713_assgn67131 <= z6713_assgn67130;
        z6713_assgn67132 <= z6713_assgn67131;
        z6713_assgn67133 <= z6713_assgn67132;
        z6713_assgn67134 <= z6713_assgn67133;
        z6713_assgn67135 <= z6713_assgn67134;
        z6713_assgn67136 <= z6713_assgn67135;
        z6713_assgn67137 <= z6713_assgn67136;
        z6713_assgn67138 <= z6713_assgn67137;
        z2651_assgn2651 <= z6713_assgn67138;
        z6725_assgn67250 <= z6725_assgn6725;
        z6725_assgn67251 <= z6725_assgn67250;
        z6725_assgn67252 <= z6725_assgn67251;
        z6725_assgn67253 <= z6725_assgn67252;
        z6725_assgn67254 <= z6725_assgn67253;
        z6725_assgn67255 <= z6725_assgn67254;
        z6725_assgn67256 <= z6725_assgn67255;
        z6725_assgn67257 <= z6725_assgn67256;
        z6725_assgn67258 <= z6725_assgn67257;
        z2661_assgn2661 <= z6725_assgn67258;
        z6729_assgn67290 <= z6729_assgn6729;
        z6729_assgn67291 <= z6729_assgn67290;
        z6729_assgn67292 <= z6729_assgn67291;
        z6729_assgn67293 <= z6729_assgn67292;
        z6729_assgn67294 <= z6729_assgn67293;
        z6729_assgn67295 <= z6729_assgn67294;
        z6729_assgn67296 <= z6729_assgn67295;
        z6729_assgn67297 <= z6729_assgn67296;
        z6729_assgn67298 <= z6729_assgn67297;
        z2663_assgn2663 <= z6729_assgn67298;
        z6737_assgn67370 <= z6737_assgn6737;
        z6737_assgn67371 <= z6737_assgn67370;
        z6737_assgn67372 <= z6737_assgn67371;
        z6737_assgn67373 <= z6737_assgn67372;
        z6737_assgn67374 <= z6737_assgn67373;
        z6737_assgn67375 <= z6737_assgn67374;
        z6737_assgn67376 <= z6737_assgn67375;
        z6737_assgn67377 <= z6737_assgn67376;
        z2669_assgn2669 <= z6737_assgn67377;
        z6741_assgn67410 <= z6741_assgn6741;
        z6741_assgn67411 <= z6741_assgn67410;
        z6741_assgn67412 <= z6741_assgn67411;
        z6741_assgn67413 <= z6741_assgn67412;
        z6741_assgn67414 <= z6741_assgn67413;
        z6741_assgn67415 <= z6741_assgn67414;
        z6741_assgn67416 <= z6741_assgn67415;
        z6741_assgn67417 <= z6741_assgn67416;
        z2671_assgn2671 <= z6741_assgn67417;
        z6749_assgn67490 <= z6749_assgn6749;
        z6749_assgn67491 <= z6749_assgn67490;
        z6749_assgn67492 <= z6749_assgn67491;
        z6749_assgn67493 <= z6749_assgn67492;
        z6749_assgn67494 <= z6749_assgn67493;
        z6749_assgn67495 <= z6749_assgn67494;
        z6749_assgn67496 <= z6749_assgn67495;
        z6749_assgn67497 <= z6749_assgn67496;
        z6749_assgn67498 <= z6749_assgn67497;
        y_G256_newbasis1 <= z6749_assgn67498;
        z6753_assgn67530 <= z6753_assgn6753;
        z6753_assgn67531 <= z6753_assgn67530;
        z6753_assgn67532 <= z6753_assgn67531;
        z6753_assgn67533 <= z6753_assgn67532;
        z6753_assgn67534 <= z6753_assgn67533;
        z6753_assgn67535 <= z6753_assgn67534;
        z6753_assgn67536 <= z6753_assgn67535;
        z6753_assgn67537 <= z6753_assgn67536;
        z6753_assgn67538 <= z6753_assgn67537;
        z2681_assgn2681 <= z6753_assgn67538;
        z6767_assgn67670 <= z6767_assgn6767;
        z6767_assgn67671 <= z6767_assgn67670;
        z6767_assgn67672 <= z6767_assgn67671;
        z6767_assgn67673 <= z6767_assgn67672;
        z6767_assgn67674 <= z6767_assgn67673;
        z6767_assgn67675 <= z6767_assgn67674;
        z6767_assgn67676 <= z6767_assgn67675;
        z6767_assgn67677 <= z6767_assgn67676;
        z6767_assgn67678 <= z6767_assgn67677;
        z2693_assgn2693 <= z6767_assgn67678;
        z6773_assgn67730 <= z6773_assgn6773;
        z6773_assgn67731 <= z6773_assgn67730;
        z6773_assgn67732 <= z6773_assgn67731;
        z6773_assgn67733 <= z6773_assgn67732;
        z6773_assgn67734 <= z6773_assgn67733;
        z6773_assgn67735 <= z6773_assgn67734;
        z6773_assgn67736 <= z6773_assgn67735;
        z6773_assgn67737 <= z6773_assgn67736;
        z6773_assgn67738 <= z6773_assgn67737;
        z2697_assgn2697 <= z6773_assgn67738;
        z6779_assgn67790 <= z6779_assgn6779;
        z6779_assgn67791 <= z6779_assgn67790;
        z6779_assgn67792 <= z6779_assgn67791;
        z6779_assgn67793 <= z6779_assgn67792;
        z6779_assgn67794 <= z6779_assgn67793;
        z6779_assgn67795 <= z6779_assgn67794;
        z6779_assgn67796 <= z6779_assgn67795;
        z6779_assgn67797 <= z6779_assgn67796;
        z6779_assgn67798 <= z6779_assgn67797;
        z2701_assgn2701 <= z6779_assgn67798;
        z6789_assgn67890 <= z6789_assgn6789;
        z6789_assgn67891 <= z6789_assgn67890;
        z6789_assgn67892 <= z6789_assgn67891;
        z6789_assgn67893 <= z6789_assgn67892;
        z6789_assgn67894 <= z6789_assgn67893;
        z6789_assgn67895 <= z6789_assgn67894;
        z6789_assgn67896 <= z6789_assgn67895;
        z6789_assgn67897 <= z6789_assgn67896;
        z6789_assgn67898 <= z6789_assgn67897;
        z2709_assgn2709 <= z6789_assgn67898;
        z6795_assgn67950 <= z6795_assgn6795;
        z6795_assgn67951 <= z6795_assgn67950;
        z6795_assgn67952 <= z6795_assgn67951;
        z6795_assgn67953 <= z6795_assgn67952;
        z6795_assgn67954 <= z6795_assgn67953;
        z6795_assgn67955 <= z6795_assgn67954;
        z6795_assgn67956 <= z6795_assgn67955;
        z6795_assgn67957 <= z6795_assgn67956;
        z6795_assgn67958 <= z6795_assgn67957;
        z2713_assgn2713 <= z6795_assgn67958;
        z6801_assgn68010 <= z6801_assgn6801;
        z6801_assgn68011 <= z6801_assgn68010;
        z6801_assgn68012 <= z6801_assgn68011;
        z6801_assgn68013 <= z6801_assgn68012;
        z6801_assgn68014 <= z6801_assgn68013;
        z6801_assgn68015 <= z6801_assgn68014;
        z6801_assgn68016 <= z6801_assgn68015;
        z6801_assgn68017 <= z6801_assgn68016;
        z2717_assgn2717 <= z6801_assgn68017;
        z6811_assgn68110 <= z6811_assgn6811;
        z6811_assgn68111 <= z6811_assgn68110;
        z6811_assgn68112 <= z6811_assgn68111;
        z6811_assgn68113 <= z6811_assgn68112;
        z6811_assgn68114 <= z6811_assgn68113;
        z6811_assgn68115 <= z6811_assgn68114;
        z6811_assgn68116 <= z6811_assgn68115;
        z6811_assgn68117 <= z6811_assgn68116;
        z6811_assgn68118 <= z6811_assgn68117;
        z2725_assgn2725 <= z6811_assgn68118;
        z6817_assgn68170 <= z6817_assgn6817;
        z6817_assgn68171 <= z6817_assgn68170;
        z6817_assgn68172 <= z6817_assgn68171;
        z6817_assgn68173 <= z6817_assgn68172;
        z6817_assgn68174 <= z6817_assgn68173;
        z6817_assgn68175 <= z6817_assgn68174;
        z6817_assgn68176 <= z6817_assgn68175;
        z6817_assgn68177 <= z6817_assgn68176;
        z6817_assgn68178 <= z6817_assgn68177;
        z2729_assgn2729 <= z6817_assgn68178;
        z6831_assgn68310 <= z6831_assgn6831;
        z6831_assgn68311 <= z6831_assgn68310;
        z6831_assgn68312 <= z6831_assgn68311;
        z6831_assgn68313 <= z6831_assgn68312;
        z6831_assgn68314 <= z6831_assgn68313;
        z6831_assgn68315 <= z6831_assgn68314;
        z6831_assgn68316 <= z6831_assgn68315;
        z6831_assgn68317 <= z6831_assgn68316;
        z6831_assgn68318 <= z6831_assgn68317;
        z2741_assgn2741 <= z6831_assgn68318;
        z6837_assgn68370 <= z6837_assgn6837;
        z6837_assgn68371 <= z6837_assgn68370;
        z6837_assgn68372 <= z6837_assgn68371;
        z6837_assgn68373 <= z6837_assgn68372;
        z6837_assgn68374 <= z6837_assgn68373;
        z6837_assgn68375 <= z6837_assgn68374;
        z6837_assgn68376 <= z6837_assgn68375;
        z6837_assgn68377 <= z6837_assgn68376;
        z6837_assgn68378 <= z6837_assgn68377;
        z2745_assgn2745 <= z6837_assgn68378;
        z6851_assgn68510 <= z6851_assgn6851;
        z6851_assgn68511 <= z6851_assgn68510;
        z6851_assgn68512 <= z6851_assgn68511;
        z6851_assgn68513 <= z6851_assgn68512;
        z6851_assgn68514 <= z6851_assgn68513;
        z6851_assgn68515 <= z6851_assgn68514;
        z6851_assgn68516 <= z6851_assgn68515;
        z6851_assgn68517 <= z6851_assgn68516;
        z6851_assgn68518 <= z6851_assgn68517;
        z2757_assgn2757 <= z6851_assgn68518;
        z6857_assgn68570 <= z6857_assgn6857;
        z6857_assgn68571 <= z6857_assgn68570;
        z6857_assgn68572 <= z6857_assgn68571;
        z6857_assgn68573 <= z6857_assgn68572;
        z6857_assgn68574 <= z6857_assgn68573;
        z6857_assgn68575 <= z6857_assgn68574;
        z6857_assgn68576 <= z6857_assgn68575;
        z6857_assgn68577 <= z6857_assgn68576;
        z6857_assgn68578 <= z6857_assgn68577;
        z2761_assgn2761 <= z6857_assgn68578;
        z6871_assgn68710 <= z6871_assgn6871;
        z6871_assgn68711 <= z6871_assgn68710;
        z6871_assgn68712 <= z6871_assgn68711;
        z6871_assgn68713 <= z6871_assgn68712;
        z6871_assgn68714 <= z6871_assgn68713;
        z6871_assgn68715 <= z6871_assgn68714;
        z6871_assgn68716 <= z6871_assgn68715;
        z6871_assgn68717 <= z6871_assgn68716;
        z6871_assgn68718 <= z6871_assgn68717;
        z2773_assgn2773 <= z6871_assgn68718;
        z6877_assgn68770 <= z6877_assgn6877;
        z6877_assgn68771 <= z6877_assgn68770;
        z6877_assgn68772 <= z6877_assgn68771;
        z6877_assgn68773 <= z6877_assgn68772;
        z6877_assgn68774 <= z6877_assgn68773;
        z6877_assgn68775 <= z6877_assgn68774;
        z6877_assgn68776 <= z6877_assgn68775;
        z6877_assgn68777 <= z6877_assgn68776;
        z6877_assgn68778 <= z6877_assgn68777;
        z2777_assgn2777 <= z6877_assgn68778;
        z6891_assgn68910 <= z6891_assgn6891;
        z6891_assgn68911 <= z6891_assgn68910;
        z6891_assgn68912 <= z6891_assgn68911;
        z6891_assgn68913 <= z6891_assgn68912;
        z6891_assgn68914 <= z6891_assgn68913;
        z6891_assgn68915 <= z6891_assgn68914;
        z6891_assgn68916 <= z6891_assgn68915;
        z6891_assgn68917 <= z6891_assgn68916;
        z6891_assgn68918 <= z6891_assgn68917;
        z2789_assgn2789 <= z6891_assgn68918;
        z6897_assgn68970 <= z6897_assgn6897;
        z6897_assgn68971 <= z6897_assgn68970;
        z6897_assgn68972 <= z6897_assgn68971;
        z6897_assgn68973 <= z6897_assgn68972;
        z6897_assgn68974 <= z6897_assgn68973;
        z6897_assgn68975 <= z6897_assgn68974;
        z6897_assgn68976 <= z6897_assgn68975;
        z6897_assgn68977 <= z6897_assgn68976;
        z6897_assgn68978 <= z6897_assgn68977;
        z2793_assgn2793 <= z6897_assgn68978;
        z6911_assgn69110 <= z6911_assgn6911;
        z6911_assgn69111 <= z6911_assgn69110;
        z6911_assgn69112 <= z6911_assgn69111;
        z6911_assgn69113 <= z6911_assgn69112;
        z6911_assgn69114 <= z6911_assgn69113;
        z6911_assgn69115 <= z6911_assgn69114;
        z6911_assgn69116 <= z6911_assgn69115;
        z6911_assgn69117 <= z6911_assgn69116;
        z6911_assgn69118 <= z6911_assgn69117;
        z2805_assgn2805 <= z6911_assgn69118;
        z6917_assgn69170 <= z6917_assgn6917;
        z6917_assgn69171 <= z6917_assgn69170;
        z6917_assgn69172 <= z6917_assgn69171;
        z6917_assgn69173 <= z6917_assgn69172;
        z6917_assgn69174 <= z6917_assgn69173;
        z6917_assgn69175 <= z6917_assgn69174;
        z6917_assgn69176 <= z6917_assgn69175;
        z6917_assgn69177 <= z6917_assgn69176;
        z6917_assgn69178 <= z6917_assgn69177;
        z_y_G256_newbasis1 <= z6917_assgn69178;
        z6921_assgn69210 <= z6921_assgn6921;
        z6921_assgn69211 <= z6921_assgn69210;
        z6921_assgn69212 <= z6921_assgn69211;
        z6921_assgn69213 <= z6921_assgn69212;
        z6921_assgn69214 <= z6921_assgn69213;
        z6921_assgn69215 <= z6921_assgn69214;
        z6921_assgn69216 <= z6921_assgn69215;
        z6921_assgn69217 <= z6921_assgn69216;
        z6921_assgn69218 <= z6921_assgn69217;
        z2813_assgn2813 <= z6921_assgn69218;
        z6935_assgn69350 <= z6935_assgn6935;
        z6935_assgn69351 <= z6935_assgn69350;
        z6935_assgn69352 <= z6935_assgn69351;
        z6935_assgn69353 <= z6935_assgn69352;
        z6935_assgn69354 <= z6935_assgn69353;
        z6935_assgn69355 <= z6935_assgn69354;
        z6935_assgn69356 <= z6935_assgn69355;
        z6935_assgn69357 <= z6935_assgn69356;
        z6935_assgn69358 <= z6935_assgn69357;
        z2825_assgn2825 <= z6935_assgn69358;
        z6941_assgn69410 <= z6941_assgn6941;
        z6941_assgn69411 <= z6941_assgn69410;
        z6941_assgn69412 <= z6941_assgn69411;
        z6941_assgn69413 <= z6941_assgn69412;
        z6941_assgn69414 <= z6941_assgn69413;
        z6941_assgn69415 <= z6941_assgn69414;
        z6941_assgn69416 <= z6941_assgn69415;
        z6941_assgn69417 <= z6941_assgn69416;
        z6941_assgn69418 <= z6941_assgn69417;
        z2829_assgn2829 <= z6941_assgn69418;
        z6947_assgn69470 <= z6947_assgn6947;
        z6947_assgn69471 <= z6947_assgn69470;
        z6947_assgn69472 <= z6947_assgn69471;
        z6947_assgn69473 <= z6947_assgn69472;
        z6947_assgn69474 <= z6947_assgn69473;
        z6947_assgn69475 <= z6947_assgn69474;
        z6947_assgn69476 <= z6947_assgn69475;
        z6947_assgn69477 <= z6947_assgn69476;
        z6947_assgn69478 <= z6947_assgn69477;
        z2833_assgn2833 <= z6947_assgn69478;
        z6957_assgn69570 <= z6957_assgn6957;
        z6957_assgn69571 <= z6957_assgn69570;
        z6957_assgn69572 <= z6957_assgn69571;
        z6957_assgn69573 <= z6957_assgn69572;
        z6957_assgn69574 <= z6957_assgn69573;
        z6957_assgn69575 <= z6957_assgn69574;
        z6957_assgn69576 <= z6957_assgn69575;
        z6957_assgn69577 <= z6957_assgn69576;
        z6957_assgn69578 <= z6957_assgn69577;
        z2841_assgn2841 <= z6957_assgn69578;
        z6963_assgn69630 <= z6963_assgn6963;
        z6963_assgn69631 <= z6963_assgn69630;
        z6963_assgn69632 <= z6963_assgn69631;
        z6963_assgn69633 <= z6963_assgn69632;
        z6963_assgn69634 <= z6963_assgn69633;
        z6963_assgn69635 <= z6963_assgn69634;
        z6963_assgn69636 <= z6963_assgn69635;
        z6963_assgn69637 <= z6963_assgn69636;
        z6963_assgn69638 <= z6963_assgn69637;
        z2845_assgn2845 <= z6963_assgn69638;
        z6969_assgn69690 <= z6969_assgn6969;
        z6969_assgn69691 <= z6969_assgn69690;
        z6969_assgn69692 <= z6969_assgn69691;
        z6969_assgn69693 <= z6969_assgn69692;
        z6969_assgn69694 <= z6969_assgn69693;
        z6969_assgn69695 <= z6969_assgn69694;
        z6969_assgn69696 <= z6969_assgn69695;
        z6969_assgn69697 <= z6969_assgn69696;
        z2849_assgn2849 <= z6969_assgn69697;
        z6979_assgn69790 <= z6979_assgn6979;
        z6979_assgn69791 <= z6979_assgn69790;
        z6979_assgn69792 <= z6979_assgn69791;
        z6979_assgn69793 <= z6979_assgn69792;
        z6979_assgn69794 <= z6979_assgn69793;
        z6979_assgn69795 <= z6979_assgn69794;
        z6979_assgn69796 <= z6979_assgn69795;
        z6979_assgn69797 <= z6979_assgn69796;
        z6979_assgn69798 <= z6979_assgn69797;
        z2857_assgn2857 <= z6979_assgn69798;
        z6985_assgn69850 <= z6985_assgn6985;
        z6985_assgn69851 <= z6985_assgn69850;
        z6985_assgn69852 <= z6985_assgn69851;
        z6985_assgn69853 <= z6985_assgn69852;
        z6985_assgn69854 <= z6985_assgn69853;
        z6985_assgn69855 <= z6985_assgn69854;
        z6985_assgn69856 <= z6985_assgn69855;
        z6985_assgn69857 <= z6985_assgn69856;
        z6985_assgn69858 <= z6985_assgn69857;
        z2861_assgn2861 <= z6985_assgn69858;
        z6999_assgn69990 <= z6999_assgn6999;
        z6999_assgn69991 <= z6999_assgn69990;
        z6999_assgn69992 <= z6999_assgn69991;
        z6999_assgn69993 <= z6999_assgn69992;
        z6999_assgn69994 <= z6999_assgn69993;
        z6999_assgn69995 <= z6999_assgn69994;
        z6999_assgn69996 <= z6999_assgn69995;
        z6999_assgn69997 <= z6999_assgn69996;
        z6999_assgn69998 <= z6999_assgn69997;
        z2873_assgn2873 <= z6999_assgn69998;
        z7005_assgn70050 <= z7005_assgn7005;
        z7005_assgn70051 <= z7005_assgn70050;
        z7005_assgn70052 <= z7005_assgn70051;
        z7005_assgn70053 <= z7005_assgn70052;
        z7005_assgn70054 <= z7005_assgn70053;
        z7005_assgn70055 <= z7005_assgn70054;
        z7005_assgn70056 <= z7005_assgn70055;
        z7005_assgn70057 <= z7005_assgn70056;
        z7005_assgn70058 <= z7005_assgn70057;
        z2877_assgn2877 <= z7005_assgn70058;
        z7019_assgn70190 <= z7019_assgn7019;
        z7019_assgn70191 <= z7019_assgn70190;
        z7019_assgn70192 <= z7019_assgn70191;
        z7019_assgn70193 <= z7019_assgn70192;
        z7019_assgn70194 <= z7019_assgn70193;
        z7019_assgn70195 <= z7019_assgn70194;
        z7019_assgn70196 <= z7019_assgn70195;
        z7019_assgn70197 <= z7019_assgn70196;
        z7019_assgn70198 <= z7019_assgn70197;
        z2889_assgn2889 <= z7019_assgn70198;
        z7025_assgn70250 <= z7025_assgn7025;
        z7025_assgn70251 <= z7025_assgn70250;
        z7025_assgn70252 <= z7025_assgn70251;
        z7025_assgn70253 <= z7025_assgn70252;
        z7025_assgn70254 <= z7025_assgn70253;
        z7025_assgn70255 <= z7025_assgn70254;
        z7025_assgn70256 <= z7025_assgn70255;
        z7025_assgn70257 <= z7025_assgn70256;
        z7025_assgn70258 <= z7025_assgn70257;
        z2893_assgn2893 <= z7025_assgn70258;
        z7039_assgn70390 <= z7039_assgn7039;
        z7039_assgn70391 <= z7039_assgn70390;
        z7039_assgn70392 <= z7039_assgn70391;
        z7039_assgn70393 <= z7039_assgn70392;
        z7039_assgn70394 <= z7039_assgn70393;
        z7039_assgn70395 <= z7039_assgn70394;
        z7039_assgn70396 <= z7039_assgn70395;
        z7039_assgn70397 <= z7039_assgn70396;
        z7039_assgn70398 <= z7039_assgn70397;
        z2905_assgn2905 <= z7039_assgn70398;
        z7045_assgn70450 <= z7045_assgn7045;
        z7045_assgn70451 <= z7045_assgn70450;
        z7045_assgn70452 <= z7045_assgn70451;
        z7045_assgn70453 <= z7045_assgn70452;
        z7045_assgn70454 <= z7045_assgn70453;
        z7045_assgn70455 <= z7045_assgn70454;
        z7045_assgn70456 <= z7045_assgn70455;
        z7045_assgn70457 <= z7045_assgn70456;
        z7045_assgn70458 <= z7045_assgn70457;
        z2909_assgn2909 <= z7045_assgn70458;
        z7059_assgn70590 <= z7059_assgn7059;
        z7059_assgn70591 <= z7059_assgn70590;
        z7059_assgn70592 <= z7059_assgn70591;
        z7059_assgn70593 <= z7059_assgn70592;
        z7059_assgn70594 <= z7059_assgn70593;
        z7059_assgn70595 <= z7059_assgn70594;
        z7059_assgn70596 <= z7059_assgn70595;
        z7059_assgn70597 <= z7059_assgn70596;
        z7059_assgn70598 <= z7059_assgn70597;
        z2921_assgn2921 <= z7059_assgn70598;
        z7065_assgn70650 <= z7065_assgn7065;
        z7065_assgn70651 <= z7065_assgn70650;
        z7065_assgn70652 <= z7065_assgn70651;
        z7065_assgn70653 <= z7065_assgn70652;
        z7065_assgn70654 <= z7065_assgn70653;
        z7065_assgn70655 <= z7065_assgn70654;
        z7065_assgn70656 <= z7065_assgn70655;
        z7065_assgn70657 <= z7065_assgn70656;
        z7065_assgn70658 <= z7065_assgn70657;
        z2925_assgn2925 <= z7065_assgn70658;
        z7079_assgn70790 <= z7079_assgn7079;
        z7079_assgn70791 <= z7079_assgn70790;
        z7079_assgn70792 <= z7079_assgn70791;
        z7079_assgn70793 <= z7079_assgn70792;
        z7079_assgn70794 <= z7079_assgn70793;
        z7079_assgn70795 <= z7079_assgn70794;
        z7079_assgn70796 <= z7079_assgn70795;
        z7079_assgn70797 <= z7079_assgn70796;
        z7079_assgn70798 <= z7079_assgn70797;
        z2937_assgn2937 <= z7079_assgn70798;
        y0 <= (t6 ^ dec_99_inp);
        y1 <= t7;
    end

endmodule

